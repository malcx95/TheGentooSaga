library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;

entity tile_and_sprite_memory is
    port (clk     : in std_logic;
          addr    : in unsigned(12 downto 0);
          pixel   : out std_logic_vector(7 downto 0);

          sprite1_addr : in unsigned(7 downto 0);
          sprite1_data : out std_logic_vector(7 downto 0));
end entity;

architecture Behavioral of tile_and_sprite_memory is
    -- Tile memory type
    type ram_t is array (0 to 8191) of std_logic_vector(7 downto 0);
    -- Sprite memory type
    type ram_s is array (0 to 1535) of std_logic_vector(7 downto 0);

    signal tile_memory : ram_t := (
            x"b1",x"8d",x"8d",x"68",x"68",x"b1",x"8d",x"8d",x"68",x"68",x"44",x"68",x"68",x"b1",x"68",x"b1",
            x"68",x"8d",x"44",x"68",x"68",x"8d",x"92",x"44",x"68",x"b1",x"8d",x"68",x"b1",x"8d",x"44",x"44",
            x"b1",x"68",x"68",x"44",x"b1",x"68",x"68",x"68",x"b1",x"68",x"68",x"68",x"44",x"44",x"b1",x"68",
            x"8d",x"6d",x"b1",x"68",x"8d",x"44",x"68",x"b1",x"8d",x"8d",x"68",x"8d",x"68",x"b1",x"8d",x"68",
            x"8d",x"68",x"8d",x"b1",x"44",x"8d",x"68",x"68",x"8d",x"44",x"68",x"6d",x"68",x"8d",x"44",x"68",
            x"68",x"44",x"8d",x"8d",x"68",x"8d",x"44",x"44",x"44",x"68",x"68",x"44",x"68",x"68",x"68",x"b1",
            x"b1",x"68",x"68",x"68",x"92",x"68",x"68",x"b1",x"b1",x"68",x"b1",x"b1",x"68",x"8d",x"68",x"8d",
            x"68",x"68",x"b1",x"b1",x"8d",x"8d",x"68",x"68",x"8d",x"44",x"8d",x"8d",x"68",x"68",x"8d",x"8d",    -- s-dirt
            x"8d",x"68",x"68",x"8d",x"68",x"8d",x"68",x"44",x"68",x"8d",x"8d",x"68",x"68",x"68",x"44",x"68",
            x"68",x"8d",x"44",x"68",x"68",x"44",x"44",x"68",x"68",x"68",x"68",x"68",x"b1",x"b1",x"68",x"8d",
            x"68",x"8d",x"68",x"b1",x"b1",x"68",x"b1",x"8d",x"44",x"b1",x"b1",x"44",x"8d",x"8d",x"92",x"68",
            x"8d",x"68",x"68",x"8d",x"8d",x"b1",x"68",x"8d",x"6d",x"8d",x"8d",x"68",x"44",x"8d",x"68",x"44",
            x"68",x"44",x"8d",x"68",x"8d",x"8d",x"b1",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"b1",x"b1",
            x"68",x"8d",x"68",x"68",x"69",x"68",x"8d",x"8d",x"68",x"44",x"b1",x"44",x"68",x"b1",x"8d",x"8d",
            x"8d",x"68",x"44",x"b1",x"68",x"44",x"68",x"44",x"b1",x"b1",x"68",x"8d",x"68",x"68",x"8d",x"8d",
            x"8d",x"68",x"b1",x"8d",x"8d",x"68",x"92",x"68",x"8d",x"8d",x"68",x"68",x"8d",x"8d",x"68",x"44",
        
            x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"54",x"50",x"50",x"50",x"50",x"50",x"2c",x"50",
            x"50",x"50",x"54",x"54",x"54",x"44",x"50",x"50",x"50",x"54",x"54",x"50",x"50",x"50",x"50",x"50",
            x"54",x"6d",x"74",x"50",x"50",x"44",x"50",x"44",x"50",x"54",x"54",x"74",x"44",x"4c",x"50",x"44",
            x"44",x"44",x"44",x"44",x"50",x"44",x"44",x"44",x"50",x"44",x"50",x"6d",x"68",x"44",x"44",x"68",
            x"68",x"44",x"8d",x"8d",x"44",x"8d",x"44",x"44",x"44",x"44",x"44",x"44",x"68",x"68",x"68",x"b1",
            x"b1",x"68",x"68",x"68",x"92",x"68",x"68",x"b1",x"b1",x"68",x"b1",x"b1",x"68",x"8d",x"68",x"8d",
            x"68",x"68",x"b1",x"b1",x"8d",x"8d",x"68",x"68",x"8d",x"44",x"8d",x"8d",x"68",x"68",x"8d",x"8d",
            x"8d",x"68",x"68",x"8d",x"68",x"8d",x"68",x"44",x"68",x"8d",x"8d",x"68",x"68",x"68",x"44",x"68",    -- s-grass
            x"68",x"8d",x"44",x"68",x"68",x"44",x"44",x"68",x"68",x"68",x"68",x"68",x"b1",x"b1",x"68",x"8d",
            x"68",x"8d",x"68",x"b1",x"b1",x"68",x"b1",x"8d",x"44",x"b1",x"b1",x"44",x"8d",x"8d",x"92",x"68",
            x"8d",x"68",x"68",x"8d",x"8d",x"b1",x"68",x"8d",x"6d",x"8d",x"8d",x"68",x"44",x"8d",x"68",x"44",
            x"68",x"44",x"8d",x"68",x"8d",x"8d",x"b1",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"b1",x"b1",
            x"68",x"8d",x"68",x"68",x"69",x"68",x"8d",x"8d",x"68",x"44",x"b1",x"44",x"68",x"b1",x"8d",x"8d",
            x"8d",x"68",x"44",x"b1",x"68",x"44",x"68",x"44",x"b1",x"b1",x"68",x"8d",x"68",x"68",x"8d",x"8d",
            x"8d",x"68",x"b1",x"8d",x"8d",x"68",x"92",x"68",x"8d",x"8d",x"68",x"68",x"8d",x"8d",x"68",x"44",
            x"68",x"68",x"68",x"8d",x"8d",x"8d",x"68",x"8d",x"68",x"92",x"92",x"44",x"68",x"8d",x"8d",x"8d",
        
            x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",
            x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",
            x"bb",x"bb",x"bb",x"db",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"df",x"bb",x"bb",x"bb",x"bb",
            x"bb",x"bb",x"db",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"df",x"bb",x"bb",x"bb",x"bb",x"bb",
            x"bb",x"df",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"df",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",
            x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"df",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",
            x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",
            x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",    -- s-ice
            x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",
            x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"df",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",
            x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"df",x"bb",x"bb",x"bb",x"bb",x"bb",x"df",x"bb",x"bb",
            x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"df",x"bb",x"bb",x"bb",
            x"bb",x"df",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"df",x"bb",x"bb",x"bb",x"bb",
            x"df",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",
            x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",
            x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",
        
            x"48",x"24",x"44",x"24",x"24",x"44",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"24",x"24",x"44",
            x"68",x"68",x"68",x"8d",x"6c",x"6c",x"8d",x"8d",x"8d",x"6c",x"48",x"44",x"44",x"48",x"68",x"68",
            x"6c",x"8d",x"48",x"24",x"24",x"44",x"44",x"24",x"24",x"44",x"68",x"68",x"68",x"68",x"68",x"68",
            x"24",x"44",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"44",x"44",x"24",x"8d",
            x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"8d",x"8d",x"8d",x"8d",x"6c",x"6c",x"68",x"24",x"24",
            x"68",x"6c",x"6c",x"8d",x"8d",x"8d",x"8d",x"44",x"24",x"68",x"68",x"6c",x"6c",x"8d",x"8d",x"68",
            x"68",x"44",x"44",x"24",x"44",x"24",x"44",x"68",x"8d",x"68",x"68",x"68",x"24",x"24",x"44",x"8d",
            x"44",x"24",x"68",x"68",x"8d",x"68",x"68",x"44",x"44",x"24",x"68",x"68",x"68",x"68",x"68",x"44",    -- s-log
            x"68",x"8d",x"68",x"24",x"24",x"24",x"68",x"68",x"8d",x"8d",x"68",x"68",x"8d",x"8d",x"8d",x"68",
            x"68",x"68",x"68",x"68",x"48",x"48",x"24",x"44",x"24",x"24",x"24",x"44",x"24",x"24",x"24",x"68",
            x"68",x"8d",x"68",x"8d",x"8d",x"8d",x"8d",x"8d",x"6c",x"6c",x"68",x"68",x"68",x"68",x"68",x"68",
            x"24",x"24",x"24",x"24",x"24",x"44",x"44",x"24",x"44",x"48",x"8d",x"8d",x"8d",x"6c",x"8d",x"6c",
            x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"24",x"24",x"24",x"24",x"44",x"44",x"68",
            x"68",x"6c",x"8d",x"68",x"8d",x"8d",x"8d",x"68",x"6c",x"6c",x"6c",x"8d",x"8d",x"6c",x"6c",x"6c",
            x"68",x"24",x"8d",x"44",x"24",x"44",x"44",x"24",x"24",x"24",x"44",x"24",x"44",x"44",x"44",x"68",
            x"6c",x"68",x"24",x"8d",x"8d",x"8d",x"6c",x"6c",x"68",x"68",x"68",x"6c",x"6c",x"8d",x"8d",x"8d",
        
            x"6d",x"ff",x"ff",x"6d",x"6d",x"ff",x"ff",x"6d",x"6d",x"ff",x"ff",x"6d",x"6d",x"ff",x"ff",x"6d",
            x"ff",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"ff",
            x"ff",x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"92",x"ff",
            x"6d",x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"92",x"6d",
            x"6d",x"92",x"ff",x"ff",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"ff",x"ff",x"92",x"6d",
            x"ff",x"92",x"ff",x"ff",x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"92",x"ff",x"ff",x"92",x"ff",
            x"ff",x"92",x"ff",x"ff",x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"92",x"ff",x"ff",x"92",x"ff",
            x"6d",x"92",x"ff",x"ff",x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"92",x"ff",x"ff",x"92",x"6d",    -- s-quartz
            x"6d",x"92",x"ff",x"ff",x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"92",x"ff",x"ff",x"92",x"6d",
            x"ff",x"92",x"ff",x"ff",x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"92",x"ff",x"ff",x"92",x"ff",
            x"ff",x"92",x"ff",x"ff",x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"92",x"ff",x"ff",x"92",x"ff",
            x"6d",x"92",x"ff",x"ff",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"ff",x"ff",x"92",x"6d",
            x"6d",x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"92",x"6d",
            x"ff",x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"92",x"ff",
            x"ff",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"ff",
            x"6d",x"ff",x"ff",x"6d",x"6d",x"ff",x"ff",x"6d",x"6d",x"ff",x"ff",x"6d",x"6d",x"ff",x"ff",x"6d",
        
            x"d6",x"fa",x"fa",x"da",x"fa",x"da",x"da",x"da",x"fa",x"da",x"da",x"da",x"da",x"ff",x"da",x"da",
            x"da",x"da",x"fa",x"fa",x"b6",x"da",x"da",x"da",x"fa",x"fa",x"ff",x"da",x"da",x"da",x"da",x"fe",
            x"fa",x"fe",x"ff",x"da",x"da",x"da",x"da",x"da",x"da",x"fa",x"fa",x"fa",x"da",x"da",x"da",x"ff",
            x"da",x"da",x"da",x"da",x"da",x"da",x"da",x"da",x"b5",x"da",x"da",x"fa",x"fa",x"fa",x"da",x"b6",
            x"fa",x"da",x"fa",x"da",x"fa",x"fa",x"fa",x"fa",x"da",x"da",x"da",x"fa",x"da",x"d6",x"fe",x"da",
            x"da",x"da",x"da",x"ff",x"da",x"fe",x"da",x"da",x"da",x"fe",x"da",x"d6",x"da",x"da",x"da",x"d6",
            x"b5",x"da",x"d6",x"da",x"b6",x"fa",x"da",x"da",x"da",x"da",x"fa",x"ff",x"da",x"fa",x"da",x"da",
            x"da",x"da",x"fa",x"da",x"da",x"da",x"fa",x"fe",x"da",x"da",x"da",x"da",x"da",x"fa",x"ff",x"fa",    -- s-sand
            x"fa",x"da",x"fe",x"fa",x"fa",x"da",x"fa",x"da",x"da",x"ff",x"d6",x"da",x"da",x"da",x"da",x"da",
            x"d6",x"da",x"fa",x"da",x"da",x"da",x"da",x"da",x"da",x"da",x"da",x"fe",x"da",x"fa",x"da",x"fe",
            x"da",x"fa",x"b5",x"fa",x"da",x"fe",x"da",x"da",x"fe",x"fe",x"fe",x"da",x"da",x"ff",x"da",x"da",
            x"da",x"fa",x"fa",x"d6",x"da",x"da",x"da",x"da",x"da",x"da",x"da",x"ff",x"da",x"da",x"da",x"b5",
            x"fe",x"da",x"da",x"fe",x"da",x"da",x"fa",x"b5",x"d6",x"da",x"da",x"da",x"fa",x"fa",x"da",x"da",
            x"da",x"fa",x"da",x"b5",x"da",x"da",x"da",x"fe",x"fa",x"fe",x"fa",x"da",x"fa",x"da",x"fa",x"da",
            x"fa",x"da",x"da",x"da",x"da",x"da",x"da",x"fa",x"da",x"da",x"b5",x"da",x"fa",x"d6",x"da",x"fa",
            x"da",x"fa",x"da",x"d6",x"ff",x"da",x"da",x"fe",x"da",x"fe",x"da",x"da",x"da",x"da",x"da",x"da",
        
            x"fa",x"fe",x"fe",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",
            x"fa",x"da",x"da",x"da",x"da",x"da",x"da",x"da",x"da",x"da",x"da",x"da",x"da",x"fa",x"fa",x"fa",
            x"da",x"da",x"da",x"d6",x"da",x"da",x"da",x"d6",x"da",x"d9",x"d5",x"d5",x"da",x"da",x"d6",x"d5",
            x"da",x"ff",x"fa",x"fe",x"d9",x"ff",x"fe",x"fe",x"fe",x"fa",x"b5",x"fe",x"fa",x"fa",x"fe",x"fe",
            x"da",x"da",x"da",x"da",x"d9",x"da",x"fa",x"fa",x"da",x"d5",x"fa",x"da",x"da",x"fa",x"da",x"da",
            x"da",x"da",x"da",x"da",x"d9",x"fa",x"da",x"fe",x"da",x"d5",x"fa",x"da",x"da",x"da",x"da",x"d5",
            x"da",x"da",x"da",x"da",x"d9",x"da",x"da",x"fa",x"b5",x"d5",x"da",x"fa",x"da",x"da",x"da",x"d5",
            x"d5",x"ff",x"fe",x"fa",x"ff",x"fe",x"da",x"da",x"fe",x"fe",x"fe",x"da",x"da",x"da",x"d5",x"fe",    -- s-sandstone
            x"fe",x"da",x"fa",x"da",x"da",x"d5",x"fe",x"fe",x"da",x"da",x"fa",x"da",x"fe",x"fe",x"d5",x"fe",
            x"da",x"fa",x"fa",x"fa",x"da",x"d5",x"fa",x"da",x"fa",x"da",x"da",x"d5",x"fa",x"da",x"d5",x"da",
            x"d5",x"d5",x"d5",x"d5",x"da",x"da",x"da",x"da",x"fa",x"da",x"da",x"da",x"da",x"d5",x"d5",x"d5",
            x"fe",x"fe",x"fe",x"fa",x"da",x"b5",x"d5",x"d5",x"da",x"d5",x"d5",x"fe",x"d5",x"fa",x"fe",x"fe",
            x"fe",x"fa",x"fa",x"da",x"fe",x"fe",x"fe",x"fe",x"d5",x"ff",x"fa",x"da",x"da",x"fa",x"fe",x"fa",
            x"fa",x"fa",x"da",x"d5",x"da",x"da",x"da",x"da",x"d5",x"da",x"da",x"da",x"d5",x"fa",x"da",x"da",
            x"da",x"da",x"fa",x"da",x"da",x"fe",x"da",x"b5",x"fa",x"d9",x"da",x"fa",x"da",x"b5",x"da",x"b5",
            x"fe",x"fe",x"da",x"da",x"da",x"da",x"d5",x"fa",x"fa",x"da",x"d5",x"da",x"fa",x"fe",x"d5",x"fe",
        
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"ff",x"ff",x"ff",x"ff",x"44",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"44",x"ff",x"ff",x"ff",x"44",x"ff",x"44",x"ff",x"ff",x"ff",x"ff",x"44",x"ff",x"ff",x"44",
            x"44",x"6d",x"44",x"44",x"ff",x"44",x"44",x"44",x"ff",x"44",x"ff",x"44",x"68",x"44",x"44",x"68",
            x"8d",x"68",x"8d",x"b1",x"44",x"8d",x"68",x"68",x"44",x"44",x"44",x"6d",x"68",x"8d",x"44",x"68",
            x"68",x"44",x"8d",x"8d",x"68",x"8d",x"44",x"44",x"44",x"68",x"68",x"44",x"68",x"68",x"68",x"b1",
            x"b1",x"44",x"68",x"68",x"92",x"68",x"68",x"b1",x"b1",x"68",x"b1",x"b1",x"68",x"8d",x"68",x"8d",
            x"b1",x"68",x"b1",x"b1",x"8d",x"8d",x"68",x"68",x"8d",x"44",x"8d",x"8d",x"68",x"68",x"8d",x"8d",    -- s-snowy-grass
            x"8d",x"68",x"68",x"8d",x"68",x"8d",x"68",x"44",x"68",x"8d",x"8d",x"68",x"68",x"68",x"44",x"68",
            x"8d",x"8d",x"44",x"68",x"68",x"44",x"44",x"68",x"68",x"68",x"68",x"68",x"b1",x"b1",x"68",x"8d",
            x"8d",x"8d",x"68",x"b1",x"b1",x"68",x"b1",x"8d",x"44",x"b1",x"b1",x"68",x"8d",x"8d",x"92",x"68",
            x"8d",x"68",x"68",x"8d",x"8d",x"b1",x"68",x"8d",x"6d",x"8d",x"8d",x"68",x"44",x"8d",x"68",x"44",
            x"68",x"44",x"8d",x"68",x"8d",x"8d",x"b1",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"b1",x"b1",
            x"68",x"8d",x"68",x"68",x"44",x"68",x"8d",x"8d",x"68",x"44",x"b1",x"44",x"68",x"b1",x"8d",x"8d",
            x"8d",x"68",x"44",x"b1",x"68",x"44",x"68",x"44",x"68",x"68",x"68",x"44",x"68",x"68",x"8d",x"8d",
            x"8d",x"68",x"b1",x"8d",x"8d",x"68",x"92",x"8d",x"8d",x"8d",x"68",x"68",x"8d",x"8d",x"68",x"44",
        
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"ff",x"ff",x"ff",x"ff",x"6d",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"6d",x"ff",x"ff",x"ff",x"6d",x"ff",x"6d",x"ff",x"ff",x"ff",x"ff",x"6d",x"ff",x"ff",x"6d",
            x"6d",x"92",x"6d",x"6d",x"ff",x"6d",x"6d",x"92",x"ff",x"6d",x"ff",x"6d",x"6d",x"6d",x"6d",x"6d",
            x"6d",x"92",x"92",x"6d",x"6d",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"6d",
            x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",
            x"92",x"92",x"6d",x"92",x"6d",x"6d",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"6d",
            x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",    -- s-snowy-stone
            x"6d",x"92",x"92",x"6d",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
            x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"6d",
            x"6d",x"6d",x"92",x"6d",x"6d",x"92",x"92",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"6d",x"6d",x"6d",
            x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"6d",x"6d",x"6d",x"92",x"92",x"6d",
            x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",
            x"6d",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",
            x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"6d",x"6d",x"6d",x"6d",
            x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",
        
            x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"6d",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",
            x"6d",x"6d",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",
            x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"6d",x"6d",
            x"6d",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",
            x"6d",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"6d",
            x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",
            x"92",x"92",x"6d",x"92",x"6d",x"6d",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"6d",
            x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",    -- s-stone
            x"6d",x"92",x"92",x"6d",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
            x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"6d",
            x"6d",x"6d",x"92",x"6d",x"6d",x"92",x"92",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"6d",x"6d",x"6d",
            x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"6d",x"6d",x"6d",x"92",x"92",x"6d",
            x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",
            x"6d",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",
            x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"6d",x"6d",x"6d",x"6d",
            x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",
        
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
        
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
        
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
        
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
        
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
        
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
            x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
        
            x"e0",x"e0",x"e0",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"bb",x"db",x"bb",x"bb",x"bb",x"bb",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"bb",x"db",x"bb",x"bb",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"bb",x"db",x"bb",x"bb",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"bb",x"db",x"bb",x"bb",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"bb",x"bb",x"bb",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"bb",x"db",x"bb",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"bb",x"bb",x"bb",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",    -- t-icicle-big
            x"e0",x"e0",x"e0",x"e0",x"e0",x"bb",x"db",x"bb",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"bb",x"db",x"bb",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"bb",x"db",x"bb",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"bb",x"db",x"bb",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"bb",x"bb",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"bb",x"bb",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"bb",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"bb",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
        
            x"e0",x"bb",x"db",x"bb",x"bb",x"bb",x"bb",x"db",x"bb",x"bb",x"bb",x"bb",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"db",x"db",x"bb",x"bb",x"e0",x"e0",x"db",x"bb",x"bb",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"bb",x"db",x"bb",x"e0",x"e0",x"e0",x"bb",x"db",x"bb",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"bb",x"db",x"bb",x"e0",x"e0",x"e0",x"bb",x"db",x"bb",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"bb",x"bb",x"bb",x"e0",x"e0",x"e0",x"e0",x"bb",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"bb",x"bb",x"e0",x"e0",x"e0",x"e0",x"bb",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"bb",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"bb",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",    -- t-icicle-small
            x"e0",x"e0",x"e0",x"bb",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
        
            x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
            x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"6d",
            x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"6d",
            x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"6d",
            x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"6d",
            x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"6d",
            x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"6d",
            x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"6d",    -- t-quartz
            x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"6d",
            x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"6d",
            x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"6d",
            x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"6d",
            x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"6d",
            x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"6d",
            x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"6d",
            x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",
        
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"14",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"14",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",    -- t-small-bush
            x"e0",x"14",x"e0",x"14",x"5d",x"e0",x"e0",x"e0",x"14",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"14",x"e0",x"14",x"e0",x"e0",x"e0",x"14",x"14",x"e0",x"e0",x"14",x"14",x"14",x"e0",x"e0",
            x"e0",x"e0",x"14",x"14",x"5d",x"e0",x"e0",x"e0",x"14",x"e0",x"e0",x"14",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"14",x"14",x"5d",x"e0",x"e0",x"14",x"e0",x"e0",x"14",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"5d",x"5d",x"14",x"14",x"14",x"14",x"5d",x"e0",x"14",x"14",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"14",x"5d",x"14",x"14",x"14",x"14",x"5d",x"e0",x"5d",x"14",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"14",x"14",x"5d",x"5d",x"14",x"14",x"14",x"14",x"14",x"5d",x"14",x"5d",x"e0",x"e0",
            x"e0",x"e0",x"14",x"14",x"5d",x"14",x"14",x"14",x"14",x"14",x"5d",x"5d",x"14",x"5d",x"e0",x"e0",
        
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",    -- t-snow
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
        
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"ff",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"ff",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",    -- t-snowy-small-bush
            x"e0",x"ff",x"e0",x"ff",x"ff",x"e0",x"e0",x"e0",x"ff",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"ff",x"e0",x"ff",x"e0",x"e0",x"e0",x"ff",x"ff",x"e0",x"e0",x"ff",x"ff",x"ff",x"e0",x"e0",
            x"e0",x"e0",x"ff",x"ff",x"5d",x"e0",x"e0",x"e0",x"ff",x"e0",x"e0",x"ff",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"ff",x"14",x"ff",x"e0",x"e0",x"ff",x"e0",x"e0",x"ff",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"ff",x"ff",x"14",x"ff",x"14",x"ff",x"ff",x"e0",x"14",x"ff",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"ff",x"5d",x"14",x"ff",x"14",x"14",x"5d",x"e0",x"5d",x"14",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"14",x"ff",x"ff",x"5d",x"14",x"14",x"ff",x"ff",x"14",x"ff",x"14",x"ff",x"e0",x"e0",
            x"e0",x"e0",x"14",x"ff",x"5d",x"14",x"14",x"14",x"14",x"14",x"ff",x"5d",x"14",x"ff",x"e0",x"e0",
        
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",    -- t-white
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
            x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
        
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
        
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
        
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
        
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
        
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
        
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
        
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
        
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
        
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
            x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0"
        );

	signal sprite_memory : ram_s := (
        x"e0",x"e0",x"e0",x"e0",x"e0",x"49",x"49",x"49",x"49",x"49",x"49",x"e0",x"e0",x"e0",x"e0",x"e0",
        x"e0",x"e0",x"e0",x"e0",x"49",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"49",x"e0",x"e0",x"e0",x"e0",
        x"e0",x"e0",x"e0",x"49",x"49",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"49",x"49",x"e0",x"e0",x"e0",
        x"e0",x"e0",x"e0",x"49",x"ff",x"ff",x"db",x"ff",x"ff",x"db",x"ff",x"b6",x"49",x"e0",x"e0",x"e0",
        x"e0",x"e0",x"e0",x"49",x"ff",x"ff",x"00",x"ff",x"ff",x"00",x"ff",x"b6",x"49",x"e0",x"e0",x"e0",
        x"e0",x"e0",x"e0",x"49",x"ff",x"ff",x"ff",x"f9",x"f9",x"ff",x"ff",x"ff",x"49",x"e0",x"e0",x"e0",
        x"e0",x"e0",x"49",x"b6",x"ff",x"ff",x"ff",x"f4",x"f4",x"ff",x"ff",x"ff",x"b6",x"49",x"e0",x"e0",
        x"e0",x"e0",x"49",x"b6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"49",x"e0",x"e0",  -- penguin
        x"e0",x"e0",x"49",x"b6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"49",x"e0",x"e0",
        x"e0",x"e0",x"49",x"b6",x"ff",x"b6",x"ff",x"ff",x"ff",x"ff",x"b6",x"ff",x"b6",x"49",x"e0",x"e0",
        x"e0",x"e0",x"49",x"b6",x"ff",x"b6",x"ff",x"ff",x"ff",x"ff",x"b6",x"ff",x"b6",x"49",x"e0",x"e0",
        x"e0",x"e0",x"49",x"49",x"b6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"49",x"49",x"e0",x"e0",
        x"e0",x"e0",x"e0",x"49",x"49",x"b6",x"ff",x"ff",x"ff",x"ff",x"b6",x"49",x"49",x"e0",x"e0",x"e0",
        x"e0",x"e0",x"e0",x"e0",x"49",x"49",x"b6",x"b6",x"b6",x"b6",x"49",x"49",x"e0",x"e0",x"e0",x"e0",
        x"e0",x"e0",x"e0",x"e0",x"f0",x"49",x"49",x"49",x"49",x"49",x"49",x"f0",x"e0",x"e0",x"e0",x"e0",
        x"e0",x"e0",x"e0",x"f0",x"f0",x"f0",x"e0",x"e0",x"e0",x"e0",x"f0",x"f0",x"f0",x"e0",x"e0",x"e0",
        
         x"e0",x"e0",x"e0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"e0",x"e0",x"e0",
         x"e0",x"e0",x"00",x"14",x"44",x"08",x"14",x"0c",x"44",x"08",x"14",x"0c",x"44",x"00",x"e0",x"e0",
         x"00",x"00",x"44",x"0c",x"0c",x"08",x"0c",x"14",x"0c",x"44",x"0c",x"08",x"0c",x"0c",x"00",x"00",
         x"00",x"0c",x"14",x"0c",x"08",x"0c",x"14",x"44",x"14",x"44",x"14",x"0c",x"44",x"14",x"0c",x"00",
         x"00",x"44",x"0c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"14",x"00",
         x"e0",x"00",x"00",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"00",x"00",x"e0",
         x"e0",x"e0",x"00",x"b6",x"b6",x"c0",x"b6",x"b6",x"b6",x"b6",x"c0",x"b6",x"b6",x"00",x"e0",x"e0",
         x"e0",x"e0",x"00",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"00",x"e0",x"e0",    -- enemy
         x"e0",x"e0",x"e0",x"00",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"00",x"e0",x"e0",x"e0",
         x"e0",x"e0",x"e0",x"e0",x"00",x"00",x"b6",x"b6",x"b6",x"b6",x"00",x"00",x"e0",x"e0",x"e0",x"e0",
         x"e0",x"00",x"e0",x"e0",x"00",x"49",x"00",x"00",x"00",x"00",x"49",x"00",x"e0",x"e0",x"00",x"e0",
         x"e0",x"e0",x"00",x"00",x"00",x"b6",x"49",x"49",x"49",x"49",x"b6",x"00",x"00",x"00",x"e0",x"e0",
         x"e0",x"00",x"e0",x"e0",x"00",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"00",x"e0",x"e0",x"00",x"e0",
         x"e0",x"e0",x"e0",x"e0",x"00",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"00",x"e0",x"e0",x"e0",x"e0",
         x"e0",x"e0",x"e0",x"e0",x"e0",x"00",x"b6",x"b6",x"b6",x"b6",x"00",x"e0",x"e0",x"e0",x"e0",x"e0",
         x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"00",x"00",x"00",x"00",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",

         x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"4a",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",
         x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"4a",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",
         x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"4a",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",
         x"e0",x"e0",x"e0",x"e0",x"e0",x"4a",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b7",
         x"e0",x"e0",x"e0",x"e0",x"4a",x"ff",x"ff",x"b7",x"b7",x"db",x"db",x"db",x"db",x"b7",x"b7",x"b7",
         x"e0",x"e0",x"e0",x"4a",x"ff",x"ff",x"93",x"b7",x"db",x"db",x"db",x"b7",x"b7",x"b7",x"b7",x"b7",
         x"e0",x"e0",x"4a",x"ff",x"ff",x"93",x"b7",x"b7",x"db",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"93",
         x"e0",x"4a",x"ff",x"ff",x"93",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"93",x"93",x"93",    -- logo-bottom-left
         x"e0",x"4a",x"ff",x"93",x"93",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"93",x"93",x"93",x"93",x"93",
         x"e0",x"4a",x"ff",x"93",x"93",x"93",x"b7",x"b7",x"b7",x"b7",x"93",x"93",x"93",x"93",x"ff",x"ff",
         x"e0",x"4a",x"ff",x"ff",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"ff",x"ff",x"ff",x"4a",
         x"e0",x"e0",x"4a",x"ff",x"ff",x"93",x"93",x"93",x"93",x"93",x"ff",x"ff",x"ff",x"4a",x"4a",x"4a",
         x"e0",x"e0",x"4a",x"4a",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"4a",x"4a",x"4a",x"e0",x"e0",
         x"e0",x"e0",x"e0",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"e0",x"e0",x"e0",x"e0",
         x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"4a",x"4a",x"4a",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
         x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",

         x"db",x"db",x"db",x"db",x"b7",x"b7",x"b7",x"93",x"93",x"93",x"93",x"ff",x"ff",x"4a",x"4a",x"e0",
         x"db",x"db",x"b7",x"b7",x"b7",x"b7",x"93",x"93",x"93",x"93",x"ff",x"ff",x"4a",x"4a",x"e0",x"e0",
         x"db",x"b7",x"b7",x"b7",x"b7",x"93",x"93",x"93",x"93",x"ff",x"ff",x"4a",x"4a",x"e0",x"e0",x"e0",
         x"b7",x"b7",x"b7",x"b7",x"93",x"93",x"93",x"93",x"ff",x"ff",x"4a",x"4a",x"e0",x"e0",x"e0",x"e0",
         x"b7",x"b7",x"b7",x"93",x"93",x"93",x"ff",x"ff",x"ff",x"4a",x"4a",x"e0",x"e0",x"e0",x"e0",x"e0",
         x"b7",x"93",x"93",x"93",x"93",x"ff",x"ff",x"4a",x"4a",x"4a",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
         x"93",x"93",x"93",x"ff",x"ff",x"ff",x"4a",x"4a",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
         x"93",x"93",x"ff",x"ff",x"4a",x"4a",x"4a",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",    -- logo-bottom-right
         x"ff",x"ff",x"ff",x"4a",x"4a",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
         x"ff",x"4a",x"4a",x"4a",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
         x"4a",x"4a",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
         x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
         x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
         x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
         x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
         x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",

         x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
         x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",
         x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"4a",x"4a",x"93",x"93",x"93",x"93",x"93",x"93",
         x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"4a",x"4a",x"93",x"93",x"93",x"93",x"b7",x"b7",x"b7",x"b7",
         x"e0",x"e0",x"e0",x"e0",x"e0",x"4a",x"4a",x"93",x"93",x"93",x"db",x"db",x"db",x"db",x"b7",x"b7",
         x"e0",x"e0",x"e0",x"e0",x"4a",x"93",x"93",x"93",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",
         x"e0",x"e0",x"e0",x"4a",x"93",x"93",x"93",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",
         x"e0",x"e0",x"4a",x"93",x"93",x"93",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"4a",    -- logo-top-left
         x"e0",x"e0",x"4a",x"93",x"93",x"93",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"4a",x"db",
         x"e0",x"4a",x"4a",x"93",x"93",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"4a",x"db",
         x"e0",x"4a",x"4a",x"93",x"93",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"4a",
         x"e0",x"e0",x"4a",x"93",x"93",x"93",x"93",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
         x"e0",x"e0",x"4a",x"4a",x"93",x"93",x"93",x"93",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
         x"e0",x"e0",x"e0",x"4a",x"4a",x"4a",x"93",x"93",x"93",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
         x"e0",x"e0",x"e0",x"e0",x"e0",x"4a",x"4a",x"4a",x"93",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",
         x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"4a",x"4a",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",

         x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
         x"4a",x"4a",x"4a",x"4a",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
         x"93",x"93",x"93",x"93",x"4a",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
         x"b7",x"b7",x"b7",x"93",x"93",x"4a",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
         x"b7",x"b7",x"b7",x"b7",x"93",x"93",x"4a",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
         x"b7",x"b7",x"b7",x"b7",x"b7",x"93",x"ff",x"4a",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
         x"db",x"db",x"b7",x"b7",x"b7",x"b7",x"93",x"ff",x"4a",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
         x"4a",x"db",x"db",x"b7",x"b7",x"b7",x"93",x"93",x"ff",x"4a",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",    -- logo-top-right
         x"db",x"4a",x"db",x"b7",x"b7",x"b7",x"b7",x"93",x"93",x"ff",x"4a",x"e0",x"e0",x"e0",x"e0",x"e0",
         x"93",x"4a",x"db",x"db",x"b7",x"b7",x"b7",x"b7",x"93",x"93",x"ff",x"4a",x"e0",x"e0",x"e0",x"e0",
         x"4a",x"ff",x"db",x"db",x"b7",x"b7",x"b7",x"b7",x"b7",x"93",x"93",x"ff",x"4a",x"e0",x"e0",x"e0",
         x"ff",x"ff",x"db",x"db",x"db",x"b7",x"b7",x"b7",x"b7",x"b7",x"93",x"93",x"ff",x"4a",x"e0",x"e0",
         x"ff",x"db",x"db",x"db",x"db",x"db",x"b7",x"b7",x"b7",x"b7",x"93",x"93",x"93",x"ff",x"4a",x"e0",
         x"db",x"db",x"db",x"db",x"db",x"db",x"b7",x"b7",x"b7",x"b7",x"93",x"93",x"93",x"ff",x"4a",x"e0",
         x"db",x"db",x"db",x"db",x"db",x"b7",x"b7",x"b7",x"b7",x"93",x"93",x"93",x"93",x"ff",x"4a",x"e0",
         x"db",x"db",x"db",x"db",x"db",x"b7",x"b7",x"b7",x"93",x"93",x"93",x"93",x"ff",x"ff",x"4a",x"e0"

    );


begin
    process(clk)
    begin
        if rising_edge(clk) then
            pixel <= tile_memory(to_integer(addr));
            sprite1_data <= sprite_memory(to_integer(sprite1_addr));
        end if;
    end process;

end Behavioral;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity pict_mem is
    port (
        clk      : in std_logic;
        data_out : out std_logic_vector(4 downto 0);
        addr    : in unsigned(11 downto 0)
        -- TODO: add sidescrolling
         );
end pict_mem;

architecture Behavioral of pict_mem is
    type ram_t is array (0 to 2249) of std_logic_vector(4 downto 0);
    signal pictMem : ram_t := (0 => "00000",1 => "00000",2 => "00000",3 => "00000",4 => "00000",5 => "00000",6 => "00000",7 => "00000",8 => "00000",9 => "00000",10 => "00000",11 => "00000",12 => "00000",13 => "00000",14 => "00000",15 => "00000",16 => "00000",17 => "00000",18 => "00000",19 => "00000",
    20 => "00000",21 => "00000",22 => "00000",23 => "00000",24 => "00000",25 => "00000",26 => "00000",27 => "00000",28 => "00001",29 => "00001",30 => "00001",31 => "00000",32 => "00000",33 => "00000",34 => "00000",35 => "00000",36 => "00000",37 => "00000",38 => "00000",39 => "00000",
    40 => "00000",41 => "00000",42 => "00000",43 => "00000",44 => "00000",45 => "00000",46 => "00000",47 => "00000",48 => "00000",49 => "00001",50 => "00000",51 => "00000",52 => "00000",53 => "00000",54 => "00000",55 => "00000",56 => "00000",57 => "00000",58 => "00000",59 => "00000",
    60 => "00000",61 => "00000",62 => "00000",63 => "00000",64 => "00000",65 => "00000",66 => "00000",67 => "00000",68 => "00000",69 => "00001",70 => "00000",71 => "00000",72 => "00000",73 => "00000",74 => "00000",75 => "00000",76 => "00000",77 => "00000",78 => "00000",79 => "00000",
    80 => "00000",81 => "00000",82 => "00000",83 => "00000",84 => "00000",85 => "00000",86 => "00000",87 => "00000",88 => "00001",89 => "00001",90 => "00001",91 => "00000",92 => "00000",93 => "00000",94 => "00000",95 => "00000",96 => "00000",97 => "00000",98 => "00000",99 => "00000",
    100 => "00000",101 => "00000",102 => "00000",103 => "00000",104 => "00000",105 => "00000",106 => "00000",107 => "00000",108 => "00000",109 => "00000",110 => "00000",111 => "00000",112 => "00000",113 => "00000",114 => "00000",115 => "00000",116 => "00000",117 => "00000",118 => "00000",119 => "00000",
    120 => "00000",121 => "00000",122 => "00010",123 => "00000",124 => "00010",125 => "00000",126 => "00010",127 => "00010",128 => "00010",129 => "00000",130 => "00010",131 => "00010",132 => "00010",133 => "00000",134 => "00010",135 => "00000",136 => "00010",137 => "00000",138 => "00000",139 => "00000",
    140 => "00000",141 => "00000",142 => "00010",143 => "00000",144 => "00010",145 => "00000",146 => "00010",147 => "00000",148 => "00010",149 => "00000",150 => "00010",151 => "00000",152 => "00000",153 => "00000",154 => "00010",155 => "00010",156 => "00000",157 => "00000",158 => "00000",159 => "00000",
    160 => "00000",161 => "00000",162 => "00010",163 => "00010",164 => "00010",165 => "00000",166 => "00010",167 => "00010",168 => "00010",169 => "00000",170 => "00010",171 => "00000",172 => "00000",173 => "00000",174 => "00010",175 => "00000",176 => "00010",177 => "00000",178 => "00000",179 => "00000",
    180 => "00000",181 => "00000",182 => "00010",183 => "00000",184 => "00010",185 => "00000",186 => "00010",187 => "00000",188 => "00010",189 => "00000",190 => "00010",191 => "00010",192 => "00010",193 => "00000",194 => "00010",195 => "00000",196 => "00010",197 => "00000",198 => "00000",199 => "00000",
    200 => "00000",201 => "00000",202 => "00000",203 => "00000",204 => "00000",205 => "00000",206 => "00000",207 => "00000",208 => "00000",209 => "00000",210 => "00000",211 => "00000",212 => "00000",213 => "00000",214 => "00000",215 => "00000",216 => "00000",217 => "00000",218 => "00000",219 => "00000",
    220 => "00000",221 => "00000",222 => "00000",223 => "00000",224 => "00001",225 => "00000",226 => "00001",227 => "00000",228 => "00001",229 => "00001",230 => "00001",231 => "00000",232 => "00001",233 => "00000",234 => "00001",235 => "00000",236 => "00000",237 => "00000",238 => "00000",239 => "00000",
    240 => "00000",241 => "00000",242 => "00000",243 => "00000",244 => "00001",245 => "00000",246 => "00001",247 => "00000",248 => "00001",249 => "00000",250 => "00001",251 => "00000",252 => "00001",253 => "00000",254 => "00001",255 => "00000",256 => "00000",257 => "00000",258 => "00000",259 => "00000",
    260 => "00000",261 => "00000",262 => "00000",263 => "00000",264 => "00000",265 => "00001",266 => "00000",267 => "00000",268 => "00001",269 => "00000",270 => "00001",271 => "00000",272 => "00001",273 => "00000",274 => "00001",275 => "00000",276 => "00000",277 => "00000",278 => "00000",279 => "00000",
    280 => "00000",281 => "00000",282 => "00000",283 => "00000",284 => "00000",285 => "00001",286 => "00000",287 => "00000",288 => "00001",289 => "00001",290 => "00001",291 => "00000",292 => "00001",293 => "00001",294 => "00001",295 => "00000",296 => "00000",297 => "00000",298 => "00000",299 => "00000", others =>(others => '0'));
begin
    process(clk)
    begin
        if rising_edge(clk) then
            data_out <= pictMem(to_integer(addr));
        end if;
    end process;
end Behavioral;

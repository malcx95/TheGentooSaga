library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;

entity background_memory is
    port (clk      : in std_logic;
          addr     : in unsigned(12 downto 0);
          pixel    : out std_logic_vector(7 downto 0);
          data_out : out std_logic_vector(4 downto 0);
          bg_picture_addr : in unsigned(11 downto 0)
      );


end entity;

architecture Behavioral of background_memory is
    type ram_b is array (0 to 1279) of std_logic_vector(7 downto 0);
    type background_type is array (0 to 2249) of std_logic_vector(4 downto 0);


    -- "tileminne"-ish
    signal background_memory : ram_b := (
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",    -- aaa-empty_sky
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",

    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"ff",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"ff",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"ff",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"ff",x"ff",x"01",x"ff",x"ff",x"01",x"01",x"01",x"01",x"01",x"01",    -- bg-star-1
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"ff",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"ff",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"ff",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",

    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"df",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"df",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"df",x"df",x"df",x"01",x"df",x"df",x"df",x"01",x"01",x"01",x"01",x"01",x"01",    -- bg-star-2
    x"01",x"01",x"01",x"01",x"01",x"01",x"df",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"df",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",

    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"ff",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",    -- bg-star-3
    x"01",x"01",x"01",x"01",x"01",x"ff",x"01",x"ff",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"ff",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",

    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"df",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"df",x"01",x"df",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"df",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",    -- bg-star-4
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"df",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"df",x"01",x"df",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"df",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01"
    );
    
    -- "levelminne"-ish
    signal background_picture : background_type := (
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00010","00000","00000",
    "00011","00000","00000","00011","00000",
    "00000","00100","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00011",
    "00000","00000","00000","00000","00000",
    "00000","00000","00010","00000","00000",
    "00000","00000","00001","00000","00000",
    "00000","00000","00001","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00011","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00001","00000",
    "00000","00000","00000","00000","00001",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00001",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00010","00000","00000",
    "00000","00000","00100","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00001","00000","00100",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00011","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00100","00000","00000","00100",
    "00100","00000","00100","00000","00000",
    "00000","00010","00000","00000","00000",
    "00000","00000","00100","00000","00000",
    "00010","00000","00010","00000","00000",
    "00000","00000","00000","00010","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00010","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00100",
    "00001","00000","00001","00000","00000",
    "00000","00011","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00010","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00100","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00001","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00011","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00010","00000","00000","00011","00000",
    "00000","00000","00000","00011","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00001","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00010","00000","00011","00000","00000",
    "00000","00000","00000","00000","00010",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00011",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00001","00000","00000",
    "00000","00000","00000","00100","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00010","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00001","00010",
    "00000","00000","00000","00000","00010",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00010","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00001","00000","00000","00000","00000",
    "00011","00000","00000","00000","00000",
    "00000","00000","00001","00000","00000",
    "00100","00000","00000","00000","00000",
    "00000","00000","00001","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00001","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00001","00000","00000","00000","00001",
    "00000","00000","00000","00000","00001",
    "00010","00000","00000","00001","00000",
    "00000","00000","00001","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00100",
    "00000","00000","00000","00000","00000",
    "00000","00000","00011","00000","00000",
    "00000","00000","00000","00000","00100",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00010","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00001","00011","00000","00001",
    "00000","00000","00000","00000","00000",
    "00100","00000","00011","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00010",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00100","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00011",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00100",
    "00000","00000","00000","00000","00010",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00001",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00001",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00100","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00001","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00010",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00001",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00011","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00011","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00100","00000","00000",
    "00000","00000","00000","00001","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00001","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00001","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00011","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00100",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00100","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00010","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00001","00000","00000","00000","00011",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00010","00000","00000","00000","00001",
    "00000","00000","00000","00000","00000",
    "00000","00010","00000","00000","00000",
    "00010","00000","00000","00010","00001",
    "00000","00011","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00100",
    "00000","00000","00000","00000","00000",
    "00010","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00100","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00001","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00100","00000","00000",
    "00000","00000","00000","00010","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00011","00000","00000",
    "00000","00000","00000","00000","00000",
    "00011","00000","00000","00000","00000",
    "00011","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00011","00010","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00100",
    "00000","00000","00000","00100","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00100","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00010",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00100","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00010","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00011","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00001","00010","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00011","00000","00001","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00011",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00001","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00011","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00011",
    "00000","00000","00000","00000","00000",
    "00011","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00011","00011",
    "00000","00000","00000","00000","00000",
    "00000","00100","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00100","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00100","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00100","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00001","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00001","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00011",
    "00000","00010","00000","00000","00000",
    "00001","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00011","00000","00010","00000","00000",
    "00000","00000","00000","00000","00100",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00011","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00001","00001","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00011",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00100",
    "00000","00000","00000","00000","00000",
    "00000","00001","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00011",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00001","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00010","00000","00011",
    "00001","00000","00000","00000","00000",
    "00001","00000","00000","00000","00000",
    "00000","00000","00000","00001","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00010","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00000","00000","00000","00000",
    "00000","00011","00000","00000","00000",
    "00000","00000","00000","00000","00000"
);


begin
    process(clk)
    begin
        if rising_edge(clk) then
            pixel <= background_memory(to_integer(addr));
            data_out <= background_picture(to_integer(bg_picture_addr));
        end if;
    end process;
end Behavioral;

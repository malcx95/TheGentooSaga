library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity level_mem is
    port (
        clk      : in std_logic;
        data_out : out std_logic_vector(4 downto 0);
        addr    : in unsigned(11 downto 0);
        query_addr : in unsigned(11 downto 0);
        query_result : out std_logic
         );
end level_mem;

architecture Behavioral of level_mem is
    type ram_t is array (0 to 2249) of std_logic_vector(4 downto 0);
    signal pictMem : ram_t := (
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 00101, 11111, 
           00101, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 10000, 11111, 
           11111, 10000, 11111, 11111, 
           11111, 00101, 11111, 11111, 
           11111, 00101, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 00100, 10000, 
           10000, 00100, 11111, 11111, 
           11111, 00101, 00101, 00101, 
           00101, 00101, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 00001, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 00100, 00100, 
           00100, 00100, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 00010, 00010, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 00001, 
           00001, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 00100, 00011, 
           00011, 00100, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 00010, 00010, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 00001, 00001, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 00100, 00011, 
           00011, 00100, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           00010, 00010, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 10000, 10000, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 00000, 
           00000, 11111, 11111, 11111, 
           11111, 10000, 10000, 11111, 
           10000, 10000, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 00100, 00011, 
           00011, 00100, 10000, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 10000, 
           10000, 11111, 11111, 11111, 
           11111, 11111, 10000, 10000, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 10000, 11111, 
           11111, 10000, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 00000, 
           00010, 11111, 11111, 11111, 
           11111, 11111, 11111, 10000, 
           10000, 11111, 11111, 11111, 
           11111, 10000, 11111, 11111, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 10000, 
           10000, 10000, 10000, 11111, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 11111, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 11111, 
           00001, 00001, 00001, 00001, 
           00010, 00010, 00010, 00010, 
           00010, 00010, 00010, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00010, 
           11111, 11111, 11111, 11111, 
           11111, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00101, 00001, 00101, 00001, 
           00101, 00101, 00101, 00101, 
           00101, 11111, 00101, 00101, 
           00101, 00001, 00001, 00011, 
           00011, 00011, 00011, 00011, 
           00011, 00011, 00011, 11111, 
           00001, 00001, 00001, 00001, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00101, 00101, 00101, 00001, 
           00001, 00001, 00001, 00001, 
           00101, 00101, 00101, 00101, 
           00101, 00101, 00101, 00101, 
           00101, 00101, 00101, 00101, 
           11111, 11111, 11111, 11111, 
           11111, 00101, 00101, 00101, 
           00101, 00101, 00101, 00101, 
           00101, 00101, 00101, 00101, 
           00101, 00101, 00101, 00101, 
           00101, 00101, 00101, 00101, 
           00101, 00101, 00101, 00101, 
           00101, 00001, 00001, 00001, 
           00101, 00101, 00101, 00101, 
           00101, 11111, 00101, 00101, 
           00101, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00011, 00011, 11111, 
           00001, 00001, 00001, 00001, 
           11111, 11111, 11111, 11111, 
           11111, 11111, 11111, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00001, 
           00001, 00001, 00001, 00101, 
           00101, 00101, 00101, 00101, 
           00101, 00101, 00101, 00101, 
           00101, 00101, 00101, 00101, 
           11111, 11111, 11111, 11111, 
           11111, 00101, 00101, 00101, 
           00101, 00101, 00101, 00101, 
           00101, 00101, 00101, 00101, 
           00101, 00101, 00101, 00101, 
           00101, 00101, 00101, 00101, 
           00101, 00101, 00101, 00101
);

signal query_help : std_logic_vector(4 downto 0);

begin
    process(clk)
    begin
        if rising_edge(clk) then
            data_out <= pictMem(to_integer(addr));
            query_help <= pictMem(to_integer(query_addr));
        end if;
    end process;

    query_result <= '0' when query_help > 15 else '1';

end Behavioral;

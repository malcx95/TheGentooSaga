
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity program_memory is
    port (clk : in std_logic;
          address : in unsigned(10 downto 0);
          data : out std_logic_vector(31 downto 0));
end program_memory;

architecture Behavioral of program_memory is
    constant nop : std_logic_vector(31 downto 0) := x"54000000";

    type memory_type is array (0 to 22) of std_logic_vector(31 downto 0);
    signal program_memory : memory_type := (
	"10011101011010110000000011100000",	-- 			ADDI    R11, R11, 224
	"10011110100101000000000000000000",	-- 			ADDI	R20, R20, GENTOO_BEGINS
	"10011110101101010000000000000001",	-- 			ADDI	R21, R21, SHIT_SONG
	"11010101000000000101100000001010",	--             SW      R0, R11, SPRITE1_Y
	"11010100111000001010011111111111",	-- 			SW		R0, R20, SONG_CHOICE
	"10000111111000000100000000001000",	-- LOOP:       LW      R31, R0, NEW_FRAME
	"10111100000111110000000000000000",	--             SFEQI   R31, 0
	"00010011111111111111111111111110",	--             BF      LOOP
	"01010100000000000000000000000000",	--             NOP
	"10000100001000001000000000000000",	--             LW      R1, R0, LEFT
	"11100001010010100000100000000000",	-- 	        ADD	    R10, R10, R1
	"10000100001000001000000000000001",	-- 	        LW      R1, R0, RIGHT
	"11100001010010100000100000000010",	-- 	        SUB	    R10, R10, R1
	"11010101000000000101000000001001",	--             SW      R0, R10, SPRITE1_X
	"10000111001000001000000000000010",	-- 			LW		R25, R0, SPACE
	"10111100001110010000000000000000",	-- 			SFNEI	R25, 0
	"00010000000000000000000000000100",	-- 			BF		SONG_CHANGE
	"01010100000000000000000000000000",	-- 			NOP
	"00000011111111111111111111110011",	-- 			JMP		LOOP
	"01010100000000000000000000000000",	-- 			NOP
	"11010100111000001010111111111111",	-- SONG_CHANGE: SW		R0, R21, SONG_CHOICE
	"00000011111111111111111111110000",	--             JMP     LOOP
	"01010100000000000000000000000000"	--             NOP
 );

begin
    process(clk)
    begin
        if (rising_edge(clk)) then
            if (address >= 4 and address <= 22) then
                data <= program_memory(to_integer(address - 4));
            else
                data <= nop;
            end if;
        end if;
    end process;
end Behavioral;

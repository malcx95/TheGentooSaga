
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity program_memory is
    port (clk : in std_logic;
          address : in unsigned(10 downto 0);
          data : out std_logic_vector(31 downto 0));
end program_memory;

architecture Behavioral of program_memory is
    constant nop : std_logic_vector(31 downto 0) := x"54000000";

    type memory_type is array (0 to 77) of std_logic_vector(31 downto 0);
    signal program_memory : memory_type := (
	"10011110100101000000000000000000",	-- 	ADDI	GENTOO_BEGINS_REG, GENTOO_BEGINS_REG, GENTOO_BEGINS
	"10011110110000000000000000000000",	-- 	ADDI	CURRENT_SONG_REG, ZERO, GENTOO_BEGINS 
	"11010100111000001010011111111111",	-- 	SW		ZERO, GENTOO_BEGINS_REG, SONG_CHOICE
	"10011100111000000000000011100000",	-- 	ADDI	GROUND_REG, ZERO, GROUND
	"11010101000000000011100000001010",	--     SW      ZERO, GROUND_REG, SPRITE1_Y
	"11010101000000000110000000001011",	--     SW      ZERO, SCROLL_OFFSET_REG, SCROLL_OFFSET
	"10000111111000000100000000001000",	-- LOOP: LW      NEW_FRAME_REG, ZERO, NEW_FRAME
	"10111100000111110000000000000000",	--     SFEQI   NEW_FRAME_REG, 0
	"00010011111111111111111111111110",	--     BF      LOOP
	"01010100000000000000000000000000",	--     NOP
	"11100000010011000101000000000000",	--     ADD ABS_POS_X, SCROLL_OFFSET_REG, SPRITE1_X_REG
	"11010101000000000001000000001100",	-- 	SW ZERO, ABS_POS_X, QUERY_X
	"11010101000000000010100000001101",	--     SW ZERO, HEIGHT, QUERY_Y
	"10000100100000000100000000001110",	--     LW QUERY_RES_REG, ZERO, QUERY_RES
	"10111100001001000000000000000000",	--     SFNEI QUERY_RES_REG, 0
	"00010000000000000000000000001010",	--     BF BLOCKED
	"10011100011001010000000000001111",	--     ADDI CORNER_CHK_Y, HEIGHT, 15
	"11010101000000000010100000001101",	--     SW ZERO, HEIGHT, QUERY_Y
	"10000100100000000100000000001110",	-- 	LW QUERY_RES_REG, ZERO, QUERY_RES
	"10111100001001000000000000000000",	--     SFNEI QUERY_RES_REG, 0
	"00010000000000000000000000000100",	-- 	BF BLOCKED
	"01010100000000000000000000000000",	--     NOP
	"00000000000000000000000000000011",	--     JMP END_OF_CAN_GO_SIDE
	"01010100000000000000000000000000",	--     NOP
	"10111100000000000000000000000000",	-- BLOCKED:    SFEQI, ZERO, 0
	"00010000000000000000000000001010",	--     BF NO_LEFT
	"01010100000000000000000000000000",	--     NOP
	"10000100001000001000000000000000",	-- 	LW      LR_BUTTONS, ZERO, LEFT
	"10111100000010100000000001010000",	-- 	SFEQI   SPRITE1_X_REG,LEFT_EDGE
	"00010000000000000000000000000101",	-- 	BF      SCROLL_LEFT
	"01010100000000000000000000000000",	-- 	NOP
	"11100001010010100000100000000000",	-- 	ADD	    SPRITE1_X_REG, SPRITE1_X_REG, LR_BUTTONS
	"00000000000000000000000000000011",	-- 	JMP     END_OF_LEFT
	"01010100000000000000000000000000",	-- 	NOP
	"11100001100011000000100000000000",	-- SCROLL_LEFT: ADD    SCROLL_OFFSET_REG, SCROLL_OFFSET_REG, LR_BUTTONS
	"10011100010000100000000000010000",	-- NO_LEFT: ADDI ABS_POS_X, ABS_POS_X, 16
	"11010101000000000001000000001100",	-- 	SW ZERO, ABS_POS_X, QUERY_X
	"11010101000000000010100000001101",	--     SW ZERO, HEIGHT, QUERY_Y
	"10000100100000000100000000001110",	--     LW QUERY_RES_REG, ZERO, QUERY_RES
	"10111100001001000000000000000000",	--     SFNEI QUERY_RES_REG, 0
	"00010000000000000000000000001010",	--     BF BLOCKED
	"10011100011001010000000000001111",	--     ADDI CORNER_CHK_Y, HEIGHT, 15
	"11010101000000000010100000001101",	--     SW ZERO, HEIGHT, QUERY_Y
	"10000100100000000100000000001110",	-- 	LW QUERY_RES_REG, ZERO, QUERY_RES
	"10111100001001000000000000000000",	--     SFNEI QUERY_RES_REG, 0
	"00010000000000000000000000000100",	-- 	BF BLOCKED
	"01010100000000000000000000000000",	--     NOP
	"00000000000000000000000000000011",	--     JMP END_OF_CAN_GO_SIDE
	"01010100000000000000000000000000",	--     NOP
	"10111100000000000000000000000000",	-- BLOCKED:    SFEQI, ZERO, 0
	"00010000000000000000000000001010",	--     BF NO_RIGHT
	"01010100000000000000000000000000",	--     NOP
	"10000100001000001000000000000001",	--     LW      LR_BUTTONS, ZERO, RIGHT
	"10111100000010100000000011110000",	-- 	SFEQI   SPRITE1_X_REG, RIGHT_EDGE
	"00010000000000000000000000000101",	-- 	BF      SCROLL_RIGHT
	"01010100000000000000000000000000",	-- 	NOP
	"11100001010010100000100000000010",	-- 	SUB	    SPRITE1_X_REG, SPRITE1_X_REG, LR_BUTTONS
	"00000000000000000000000000000011",	-- 	JMP     END_OF_RIGHT
	"01010100000000000000000000000000",	-- 	NOP
	"11100001100011000000100000000010",	-- SCROLL_RIGHT: SUB    SCROLL_OFFSET_REG, SCROLL_OFFSET_REG, LR_BUTTONS
	"11010101000000000101000000001001",	-- NO_RIGHT:   SW      ZERO, SPRITE1_X_REG, SPRITE1_X
	"11010101000000000110000000001011",	-- 	SW      ZERO, SCROLL_OFFSET_REG, SCROLL_OFFSET
	"10000111001000001000000000000010",	-- 	LW		SPACE_REG, ZERO, SPACE
	"11010101000000001100100000000000",	-- 	SW		ZERO, SPACE_REG, LED0
	"11100100011001110010100000000000",	-- 	SFGEU	GROUND_REG, HEIGHT
	"00010000000000000000000000001001",	-- 	BF		OFF_GROUND
	"01010100000000000000000000000000",	-- 	NOP
	"00011000101000000000000000000000",	-- 	MOVHI	HEIGHT, 0
	"11100000101000000011100000000000",	-- 	ADD		HEIGHT, ZERO, GROUND_REG
	"00011000110000000000000000000000",	-- 	MOVHI	SPEED, 0
	"10111100000110010000000000000000",	-- 	SFEQI	SPACE_REG, 0
	"00010000000000000000000000000100",	-- 	BF		NO_JUMP
	"01010100000000000000000000000000",	-- 	NOP
	"10011100110000000000000000001100",	-- 	ADDI	SPEED, ZERO, V0
	"10010100110001100000000000000001",	-- OFF_GROUND:		SUBI	SPEED, SPEED, G
	"11100000101001010011000000000010",	-- NO_JUMP:		SUB		HEIGHT, HEIGHT, SPEED
	"11010101000000000010100000001010",	-- 	SW		ZERO, HEIGHT, SPRITE1_Y
	"00000011111111111111111110111001"	-- 	JMP		LOOP
 );

begin
    process(clk)
    begin
        if (rising_edge(clk)) then
            if (address >= 4 and address <= 81) then
                data <= program_memory(to_integer(address - 4));
            else
                data <= nop;
            end if;
        end if;
    end process;
end Behavioral;

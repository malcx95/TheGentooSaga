
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity program_memory is
    port (clk : in std_logic;
          address : in unsigned(10 downto 0);
          data : out std_logic_vector(31 downto 0));
end program_memory;

architecture Behavioral of program_memory is
    constant nop : std_logic_vector(31 downto 0) := x"54000000";

    type memory_type is array (0 to 56) of std_logic_vector(31 downto 0);
    signal program_memory : memory_type := (
	"10011101011010110000000011100000",	-- 			ADDI    R11, R11, 224
	"10011110100101000000000000000000",	-- 			ADDI	R20, R20, GENTOO_BEGINS
	"10011110101101010000000000000001",	-- 			ADDI	R21, R21, SHIT_SONG
	"11100010110101000000000000000000",	-- 			ADD		R22, R20, R0 
	"11010101000000000101100000001010",	--             SW      R0, R11, SPRITE1_Y
	"11010100111000001010011111111111",	-- 			SW		R0, R20, SONG_CHOICE
	"11010101000000000110000000001011",	--             SW      R0, R12, SCROLL_OFFSET
	"10000111111000000100000000001000",	-- LOOP:       LW      R31, R0, NEW_FRAME
	"10111100000111110000000000000000",	--             SFEQI   R31, 0
	"00010011111111111111111111111110",	--             BF      LOOP
	"01010100000000000000000000000000",	--             NOP
	"10000100001000001000000000000000",	--     LW      R1, R0, LEFT
	"10111100000010100000000001010000",	--     SFEQI   R10,LEFT_EDGE
	"00010000000000000000000000000101",	--     BF      SCROLL_LEFT
	"01010100000000000000000000000000",	--     NOP
	"11100001010010100000100000000000",	-- 	ADD	    R10, R10, R1
	"00000000000000000000000000000011",	--     JMP     END_OF_LEFT
	"01010100000000000000000000000000",	--     NOP
	"11100001100011000000100000000000",	-- SCROLL_LEFT: ADD    R12, R12, R1
	"10000100001000001000000000000001",	-- END_OF_LEFT: LW      R1, R0, RIGHT
	"10111100000010100000000011110000",	--     SFEQI   R10, RIGHT_EDGE
	"00010000000000000000000000000101",	--     BF      SCROLL_RIGHT
	"01010100000000000000000000000000",	--     NOP     
	"11100001010010100000100000000010",	--     SUB	    R10, R10, R1
	"00000000000000000000000000000011",	--     JMP     END_OF_RIGHT
	"01010100000000000000000000000000",	--     NOP
	"11100001100011000000100000000010",	-- SCROLL_RIGHT: SUB    R12, R12, R1
	"11010101000000000101000000001001",	-- END_OF_RIGHT: SW      R0, R10, SPRITE1_X
	"11010101000000000110000000001011",	--     SW      R0, R12, SCROLL_OFFSET
	"10000111001000001000000000000010",	-- 			LW		R25, R0, SPACE
	"11010101000000001100100000000000",	-- 			SW		R0, R25, LED0
	"10111100001110010000000000000000",	-- 			SFNEI	R25, 0
	"00010000000000000000000000000100",	-- 			BF		SONG_CHANGE
	"01010100000000000000000000000000",	-- 			NOP
	"00000011111111111111111111100101",	-- 			JMP		LOOP
	"01010100000000000000000000000000",	-- 			NOP
	"10111100000101100000000000000000",	-- 			SFEQI	R22, GENTOO_BEGINS
	"00010000000000000000000000000101",	-- 			BF		SHIT
	"01010100000000000000000000000000",	-- 			NOP
	"00011010110000000000000000000000",	-- 			MOVHI	R22, GENTOO_BEGINS
	"00000000000000000000000000000011",	-- 			JMP		E
	"01010100000000000000000000000000",	-- 			NOP
	"10011110110000000000000000000001",	-- SHIT:		ADDI	R22, R0, SHIT_SONG
	"11010100111000001011011111111111",	-- E:			SW		R0, R22, SONG_CHOICE
	"10111100000010110000000011010110",	-- JUMP_LOOP: SFEQI   R11,214
	"00010000000000000000000000000100",	--     BF      FALL_DOWN
	"01010100000000000000000000000000",	--     NOP
	"10010101011010110000000000000001",	--     SUBI     R11,R11,1
	"00000011111111111111111111111100",	--     JMP     JUMP_LOOP
	"10111100000010110000000011100000",	-- FALL_DOWN: SFEQI   R11,224
	"00010000000000000000000000000100",	--     BF      END_JUMP
	"01010100000000000000000000000000",	--     NOP
	"10011101011010110000000000000001",	--     ADDI     R11,R11,1
	"00000011111111111111111111111101",	--     JMP    FALL_DOWN
	"01010100000000000000000000000000",	-- END_JUMP: NOP
	"00000011111111111111111111010000",	-- 			JMP		LOOP
	"01010100000000000000000000000000"	-- 			NOP
 );

begin
    process(clk)
    begin
        if (rising_edge(clk)) then
            if (address >= 4 and address <= 60) then
                data <= program_memory(to_integer(address - 4));
            else
                data <= nop;
            end if;
        end if;
    end process;
end Behavioral;

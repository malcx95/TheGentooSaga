library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;

entity music_memory is
    port (clk : in std_logic;
          address : in unsigned(6 downto 0);
          data : out unsigned(7 downto 0);
		  song_choice : in std_logic_vector(1 downto 0));

end music_memory;

architecture Behavioral of music_memory is

    type gentoo_begins_t is array (0 to 127) of unsigned(7 downto 0);

    signal gentoo_begins : gentoo_begins_t := (
        x"67", x"5f", x"58", x"66", x"58", x"5f", x"64", x"5f",
        x"6b", x"5b", x"54", x"69", x"54", x"5b", x"67", x"5b",
        x"66", x"5d", x"56", x"5d", x"56", x"5d", x"62", x"5d",
        x"5f", x"5a", x"53", x"5a", x"53", x"5a", x"53", x"5a",
        x"67", x"5f", x"58", x"66", x"58", x"5f", x"64", x"5f",
        x"6b", x"5b", x"54", x"69", x"54", x"5b", x"67", x"5b",
        x"66", x"5d", x"56", x"5d", x"56", x"5d", x"62", x"5d",
        x"5f", x"5a", x"53", x"5a", x"53", x"5a", x"53", x"5a",
        x"6b", x"5f", x"58", x"69", x"58", x"5f", x"67", x"5f",
        x"6c", x"64", x"5d", x"6b", x"5d", x"64", x"69", x"64",
        x"67", x"62", x"5b", x"69", x"5b", x"62", x"6b", x"62",
        x"66", x"5a", x"53", x"5a", x"53", x"5a", x"53", x"5a",
        x"6b", x"5f", x"58", x"69", x"58", x"5f", x"67", x"5f",
        x"6c", x"64", x"5d", x"6b", x"5d", x"64", x"69", x"64",
        x"67", x"62", x"5b", x"69", x"5b", x"62", x"6b", x"62",
        x"66", x"5a", x"53", x"5a", x"53", x"5a", x"53", x"5a");

	type example_t is array (0 to 127) of unsigned(7 downto 0);

signal example : example_t := (
"11101111", 
"11101111", "01110101", "00111101", "11100001", "00111001", "10010010", "10110101", "10001101", 
"10010100", "11011111", "01001000", "10110001", "01000010", "11011011", "10001111", "01110110", 
"11100100", "11000011", "01111101", "01101001", "10101011", "01010110", "11011011", "11001100", 
"00101110", "01110011", "00000101", "10111001", "00010011", "10001100", "00110010", "10100011", 
"00110010", "00000100", "00100011", "11111010", "00101000", "01010101", "00101111", "00101011", 
"00010001", "00001111", "10001001", "00000011", "11011101", "00100100", "00110000", "11101110", 
"10010110", "01001000", "01111000", "00100110", "10111100", "11010000", "11000011", "11000000", 
"00010011", "11000100", "00111011", "00001101", "11111111", "11101000", "10010110", "10101010", 
"10100010", "10111011", "10001101", "10110101", "01010111", "00101101", "01111110", "11010010", 
"11011100", "00101111", "00111000", "11110101", "11000010", "00000110", "10110000", "11010011", 
"10000000", "01001010", "00001110", "00010100", "00000111", "01101111", "00001010", "11100000", 
"01010010", "01100110", "10011001", "01110000", "11110110", "10111010", "11110110", "10010000", 
"10111011", "10001110", "11000011", "00011100", "10001011", "10100001", "00110010", "00001101", 
"00110010", "01011010", "01101001", "00101011", "01111110", "00001101", "01010011", "10111101", 
"10001001", "11010111", "00001011", "00000000", "00111001", "00110110", "00101010", "01011100", 
"10111001", "01000111", "10011101", "11101000", "11111110", "11110010", "11010010");

	signal song1 : unsigned(7 downto 0);
	signal song2 : unsigned(7 downto 0);

begin
    process(clk)
    begin
        if (rising_edge(clk)) then
			song1 <= gentoo_begins(to_integer(address));
			song2 <= example(to_integer(address));
        end if;
    end process;

	with song_choice select data <= 
			song1 when "00",
			song2 when "01",
			(others => '0') when others;

end Behavioral;


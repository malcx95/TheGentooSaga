
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity program_memory is
    port (clk : in std_logic;
          address : in unsigned(10 downto 0);
          data : out std_logic_vector(31 downto 0));
end program_memory;

architecture Behavioral of program_memory is
    constant nop : std_logic_vector(31 downto 0) := x"54000000";

    type memory_type is array (0 to 98) of std_logic_vector(31 downto 0);
    signal program_memory : memory_type := (
	x"9E940000",	-- 	ADDI	GENTOO_BEGINS_REG, GENTOO_BEGINS_REG, GENTOO_BEGINS
	x"9EC00000",	-- 	ADDI	CURRENT_SONG_REG, ZERO, GENTOO_BEGINS 
	x"D4E0A7FF",	-- 	SW		ZERO, GENTOO_BEGINS_REG, SONG_CHOICE
	x"9CE000A0",	-- 	ADDI	GROUND_REG, ZERO, GROUND
	x"D500380A",	--     SW      ZERO, GROUND_REG, SPRITE1_Y
	x"D500600B",	--     SW      ZERO, SCROLL_OFFSET_REG, SCROLL_OFFSET
	x"87E04008",	-- LOOP: LW      NEW_FRAME_REG, ZERO, NEW_FRAME
	x"BC1F0000",	--     SFEQI   NEW_FRAME_REG, 0
	x"13FFFFFE",	--     BF      LOOP
	x"54000000",	--     NOP
	x"E04C5000",	--     ADD ABS_POS_X, SCROLL_OFFSET_REG, SPRITE1_X_REG
	x"D500100C",	-- 	SW ZERO, ABS_POS_X, QUERY_X
	x"BC200000",	-- 	SFNEI	ZERO, 0
	x"D500280D",	--     SW ZERO, HEIGHT, QUERY_Y
	x"8480400E",	--     LW QUERY_RES_REG, ZERO, QUERY_RES
	x"BC240000",	--     SFNEI QUERY_RES_REG, 0
	x"1000000A",	--     BF XBLOCKED
	x"9C65000F",	--     ADDI CORNER_CHK_Y, HEIGHT, 15
	x"D500280D",	--     SW ZERO, HEIGHT, QUERY_Y
	x"8480400E",	-- 	LW QUERY_RES_REG, ZERO, QUERY_RES
	x"BC240000",	--     SFNEI QUERY_RES_REG, 0
	x"10000004",	-- 	BF XBLOCKED
	x"54000000",	--     NOP
	x"00000003",	--     JMP END_OF_CAN_GO_SIDE
	x"54000000",	--     NOP
	x"BC000000",	-- XBLOCKED: SFEQI, ZERO, 0
	x"1000000A",	--     BF NO_LEFT
	x"54000000",	--     NOP
	x"84208000",	-- 	LW      LR_BUTTONS, ZERO, LEFT
	x"BC0A0050",	-- 	SFEQI   SPRITE1_X_REG,LEFT_EDGE
	x"10000005",	-- 	BF      SCROLL_LEFT
	x"54000000",	-- 	NOP
	x"E14A0800",	-- 	ADD	    SPRITE1_X_REG, SPRITE1_X_REG, LR_BUTTONS
	x"00000003",	-- 	JMP     END_OF_LEFT
	x"54000000",	-- 	NOP
	x"E18C0800",	-- SCROLL_LEFT: ADD    SCROLL_OFFSET_REG, SCROLL_OFFSET_REG, LR_BUTTONS
	x"9C420010",	-- NO_LEFT: ADDI ABS_POS_X, ABS_POS_X, 16
	x"D500100C",	-- 	SW ZERO, ABS_POS_X, QUERY_X
	x"BC200000",	-- 	SFNEI	ZERO, 0
	x"D500280D",	--     SW ZERO, HEIGHT, QUERY_Y
	x"8480400E",	--     LW QUERY_RES_REG, ZERO, QUERY_RES
	x"BC240000",	--     SFNEI QUERY_RES_REG, 0
	x"1000000A",	--     BF XBLOCKED
	x"9C65000F",	--     ADDI CORNER_CHK_Y, HEIGHT, 15
	x"D500280D",	--     SW ZERO, HEIGHT, QUERY_Y
	x"8480400E",	-- 	LW QUERY_RES_REG, ZERO, QUERY_RES
	x"BC240000",	--     SFNEI QUERY_RES_REG, 0
	x"10000004",	-- 	BF XBLOCKED
	x"54000000",	--     NOP
	x"00000003",	--     JMP END_OF_CAN_GO_SIDE
	x"54000000",	--     NOP
	x"BC000000",	-- XBLOCKED: SFEQI, ZERO, 0
	x"1000000A",	--     BF NO_RIGHT
	x"54000000",	--     NOP
	x"84208001",	--     LW      LR_BUTTONS, ZERO, RIGHT
	x"BC0A00F0",	-- 	SFEQI   SPRITE1_X_REG, RIGHT_EDGE
	x"10000005",	-- 	BF      SCROLL_RIGHT
	x"54000000",	-- 	NOP
	x"E14A0802",	-- 	SUB	    SPRITE1_X_REG, SPRITE1_X_REG, LR_BUTTONS
	x"00000003",	-- 	JMP     END_OF_RIGHT
	x"54000000",	-- 	NOP
	x"E18C0802",	-- SCROLL_RIGHT: SUB    SCROLL_OFFSET_REG, SCROLL_OFFSET_REG, LR_BUTTONS
	x"D5005009",	-- NO_RIGHT:   SW      ZERO, SPRITE1_X_REG, SPRITE1_X
	x"D500600B",	-- 	SW      ZERO, SCROLL_OFFSET_REG, SCROLL_OFFSET
	x"87208002",	-- 	LW		SPACE_REG, ZERO, SPACE
	x"D500C800",	-- 	SW		ZERO, SPACE_REG, LED0
	x"9C650010",	--     ADDI    CORNER_CHK_Y, HEIGHT, 16
	x"D500180D",	--     SW      ZERO, CORNER_CHK_Y, QUERY_Y
	x"BC200000",	-- 	SFNEI	ZERO, 0
	x"E04C5000",	--     ADD ABS_POS_X, SCROLL_OFFSET_REG, SPRITE1_X_REG
	x"D500100C",	--     SW ZERO, ABS_POS_X, QUERY_X
	x"8480400E",	--     LW QUERY_RES_REG, ZERO, QUERY_RES
	x"BC240000",	--     SFNEI QUERY_RES_REG, 0
	x"10000009",	--     BF YBLOCKED
	x"9C420010",	--     ADDI ABS_POS_X, ABS_POS_X, 16
	x"D500100C",	--     SW ZERO, ABS_POS_X, QUERY_X
	x"8480400E",	--     LW QUERY_RES_REG, ZERO, QUERY_RES
	x"BC240000",	--     SFNEI QUERY_RES_REG, 0
	x"10000003",	--     BF YBLOCKED
	x"54000000",	--     NOP
	x"00000003",	--     JMP END_OF_CAN_GO_UP
	x"54000000",	--     NOP
	x"BC000000",	-- YBLOCKED: SFEQI, ZERO, 0
	x"10000005",	-- 	BF		ON_GROUND
	x"54000000",	-- 	NOP
	x"94C60001",	-- 	SUBI	SPEED, SPEED, G
	x"0000000B",	--     JMP     NO_JUMP
	x"54000000",	--     NOP
	x"54000000",	-- ON_GROUND: NOP
	x"B4A50024",	--     SRLI    HEIGHT, HEIGHT, 4
	x"B4A50004",	--     SLLI    HEIGHT, HEIGHT, 4
	x"18C00000",	-- 	MOVHI	SPEED, 0
	x"BC190000",	-- 	SFEQI	SPACE_REG, 0
	x"10000002",	-- 	BF		NO_JUMP
	x"54000000",	-- 	NOP
	x"9CC0000C",	-- 	ADDI	SPEED, ZERO, V0
	x"E0A53002",	-- NO_JUMP:		SUB		HEIGHT, HEIGHT, SPEED
	x"D500280A",	-- 	SW		ZERO, HEIGHT, SPRITE1_Y
	x"03FFFFA4"		-- 	JMP		LOOP
 );

begin
    process(clk)
    begin
        if (rising_edge(clk)) then
            if (address >= 4 and address <= 102) then
                data <= program_memory(to_integer(address - 4));
            else
                data <= nop;
            end if;
        end if;
    end process;
end Behavioral;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity level_mem is
    port (
        clk      : in std_logic;
        data_out : out std_logic_vector(4 downto 0);
        addr    : in unsigned(11 downto 0);
		query_addr : in unsigned(11 downto 0);
		query_result : out std_logic
         );
end level_mem;

architecture Behavioral of level_mem is
    type ram_t is array (0 to 2249) of std_logic_vector(4 downto 0);
    signal pictMem : ram_t := (
0=>"00000", 1=>"00000", 2=>"00000", 3=>"00000", 4=>"00000", 
5=>"00000", 6=>"00000", 7=>"00000", 8=>"00000", 9=>"00000", 
10=>"00000", 11=>"00000", 12=>"00000", 13=>"00000", 14=>"00000", 
15=>"00000", 16=>"00000", 17=>"00000", 18=>"00000", 19=>"00000", 
20=>"00000", 21=>"00000", 22=>"00000", 23=>"00000", 24=>"00000", 
25=>"00000", 26=>"00000", 27=>"00000", 28=>"00000", 29=>"00000", 
30=>"00000", 31=>"00000", 32=>"00000", 33=>"00000", 34=>"00000", 
35=>"00000", 36=>"00010", 37=>"00010", 38=>"00010", 39=>"00010", 
40=>"00000", 41=>"00000", 42=>"00000", 43=>"00000", 44=>"00000", 
45=>"00000", 46=>"00000", 47=>"00000", 48=>"00000", 49=>"00000", 
50=>"00000", 51=>"00000", 52=>"00000", 53=>"00010", 54=>"00000", 
55=>"00000", 56=>"00000", 57=>"00000", 58=>"00000", 59=>"00000", 
60=>"00000", 61=>"00000", 62=>"00000", 63=>"00000", 64=>"00000", 
65=>"00000", 66=>"00010", 67=>"00010", 68=>"00010", 69=>"00010", 
70=>"00000", 71=>"00001", 72=>"00001", 73=>"00000", 74=>"00000", 
75=>"00000", 76=>"00000", 77=>"00000", 78=>"00000", 79=>"00000", 
80=>"00000", 81=>"00000", 82=>"00000", 83=>"00000", 84=>"00000", 
85=>"00000", 86=>"00000", 87=>"00000", 88=>"00001", 89=>"00001", 
90=>"00000", 91=>"00000", 92=>"00000", 93=>"00000", 94=>"00000", 
95=>"00000", 96=>"00010", 97=>"00010", 98=>"00010", 99=>"00010", 
100=>"00000", 101=>"00001", 102=>"00001", 103=>"00000", 104=>"00000", 
105=>"00000", 106=>"00000", 107=>"00000", 108=>"00000", 109=>"00000", 
110=>"00000", 111=>"00010", 112=>"00000", 113=>"00010", 114=>"00000", 
115=>"00000", 116=>"00000", 117=>"00000", 118=>"00000", 119=>"00000", 
120=>"00000", 121=>"00001", 122=>"00000", 123=>"00000", 124=>"00001", 
125=>"00000", 126=>"00010", 127=>"00010", 128=>"00010", 129=>"00010", 
130=>"00000", 131=>"00001", 132=>"00001", 133=>"00001", 134=>"00001", 
135=>"00000", 136=>"00001", 137=>"00001", 138=>"00001", 139=>"00001", 
140=>"00000", 141=>"00000", 142=>"00000", 143=>"00000", 144=>"00000", 
145=>"00000", 146=>"00001", 147=>"00000", 148=>"00000", 149=>"00001", 
150=>"00000", 151=>"00001", 152=>"00000", 153=>"00000", 154=>"00001", 
155=>"00000", 156=>"00010", 157=>"00010", 158=>"00010", 159=>"00010", 
160=>"00000", 161=>"00001", 162=>"00001", 163=>"00001", 164=>"00001", 
165=>"00000", 166=>"00000", 167=>"00000", 168=>"00000", 169=>"00000", 
170=>"00000", 171=>"00010", 172=>"00000", 173=>"00000", 174=>"00010", 
175=>"00000", 176=>"00000", 177=>"00000", 178=>"00000", 179=>"00000", 
180=>"00000", 181=>"00000", 182=>"00000", 183=>"00000", 184=>"00000", 
185=>"00000", 186=>"00010", 187=>"00000", 188=>"00000", 189=>"00010", 
190=>"00000", 191=>"00001", 192=>"00001", 193=>"00001", 194=>"00001", 
195=>"00000", 196=>"00000", 197=>"00000", 198=>"00000", 199=>"00000", 
200=>"00000", 201=>"00000", 202=>"00000", 203=>"00000", 204=>"00000", 
205=>"00000", 206=>"00000", 207=>"00000", 208=>"00000", 209=>"00001", 
210=>"00000", 211=>"00000", 212=>"00000", 213=>"00000", 214=>"00000", 
215=>"00000", 216=>"00010", 217=>"00010", 218=>"00010", 219=>"00010", 
220=>"00000", 221=>"00001", 222=>"00001", 223=>"00001", 224=>"00001", 
225=>"00000", 226=>"00000", 227=>"00000", 228=>"00000", 229=>"00000", 
230=>"00000", 231=>"00000", 232=>"00010", 233=>"00000", 234=>"00000", 
235=>"00000", 236=>"00000", 237=>"00000", 238=>"00000", 239=>"00000", 
240=>"00000", 241=>"00000", 242=>"00000", 243=>"00000", 244=>"00000", 
245=>"00000", 246=>"00010", 247=>"00000", 248=>"00010", 249=>"00010", 
250=>"00000", 251=>"00000", 252=>"00000", 253=>"00000", 254=>"00000", 
255=>"00000", 256=>"00000", 257=>"00000", 258=>"00000", 259=>"00000", 
260=>"00000", 261=>"00000", 262=>"00000", 263=>"00000", 264=>"00000", 
265=>"00000", 266=>"00000", 267=>"00000", 268=>"00000", 269=>"00000", 
270=>"00000", 271=>"00000", 272=>"00000", 273=>"00000", 274=>"00000", 
275=>"00000", 276=>"00000", 277=>"00000", 278=>"00000", 279=>"00000", 
280=>"00000", 281=>"00000", 282=>"00000", 283=>"00000", 284=>"00000", 
285=>"00000", 286=>"00000", 287=>"00000", 288=>"00000", 289=>"00000", 
290=>"00000", 291=>"00000", 292=>"00000", 293=>"00000", 294=>"00000", 
295=>"00000", 296=>"00000", 297=>"00000", 298=>"00000", 299=>"00000", 
300=>"00101", 301=>"00101", 302=>"00101", 303=>"00101", 304=>"00101", 
305=>"00101", 306=>"00101", 307=>"00101", 308=>"00101", 309=>"00101", 
310=>"00101", 311=>"00101", 312=>"00101", 313=>"00101", 314=>"00101", 
315=>"00101", 316=>"00101", 317=>"00101", 318=>"00101", 319=>"00101", 
320=>"00101", 321=>"00101", 322=>"00101", 323=>"00101", 324=>"00101", 
325=>"00101", 326=>"00101", 327=>"00101", 328=>"00101", 329=>"00101", 
330=>"00101", 331=>"00101", 332=>"00101", 333=>"00101", 334=>"00101", 
335=>"00101", 336=>"00101", 337=>"00101", 338=>"00101", 339=>"00101", 
340=>"00101", 341=>"00101", 342=>"00101", 343=>"00101", 344=>"00101", 
345=>"00101", 346=>"00101", 347=>"00101", 348=>"00101", 349=>"00101", 
350=>"00101", 351=>"00101", 352=>"00101", 353=>"00101", 354=>"00101", 
355=>"00101", 356=>"00101", 357=>"00101", 358=>"00101", 359=>"00101", 
360=>"00101", 361=>"00101", 362=>"00101", 363=>"00101", 364=>"00101", 
365=>"00101", 366=>"00101", 367=>"00101", 368=>"00101", 369=>"00101", 
370=>"00101", 371=>"00101", 372=>"00101", 373=>"00101", 374=>"00101", 
375=>"00101", 376=>"00101", 377=>"00101", 378=>"00101", 379=>"00101", 
380=>"00101", 381=>"00101", 382=>"00101", 383=>"00101", 384=>"00101", 
385=>"00101", 386=>"00101", 387=>"00101", 388=>"00101", 389=>"00101", 
390=>"00101", 391=>"00101", 392=>"00101", 393=>"00101", 394=>"00101", 
395=>"00101", 396=>"00101", 397=>"00101", 398=>"00101", 399=>"00101", 
400=>"00101", 401=>"00101", 402=>"00101", 403=>"00101", 404=>"00101", 
405=>"00101", 406=>"00101", 407=>"00101", 408=>"00101", 409=>"00101", 
410=>"00101", 411=>"00101", 412=>"00101", 413=>"00101", 414=>"00101", 
415=>"00101", 416=>"00101", 417=>"00101", 418=>"00101", 419=>"00101", 
420=>"00101", 421=>"00101", 422=>"00101", 423=>"00101", 424=>"00101", 
425=>"00101", 426=>"00101", 427=>"00101", 428=>"00101", 429=>"00101", 
430=>"00101", 431=>"00101", 432=>"00101", 433=>"00101", 434=>"00101", 
435=>"00101", 436=>"00101", 437=>"00101", 438=>"00101", 439=>"01000", 
440=>"00101", 441=>"00101", 442=>"00101", 443=>"00101", 444=>"00101", 
445=>"00101", 446=>"00101", 447=>"00101", 448=>"00101", 449=>"00101", 
450=>"00101", 451=>"00101", 452=>"00101", 453=>"01000", 454=>"00101", 
455=>"00101", 456=>"00101", 457=>"00101", 458=>"00101", 459=>"00101", 
460=>"00101", 461=>"00101", 462=>"00101", 463=>"00101", 464=>"00101", 
465=>"00101", 466=>"01000", 467=>"01000", 468=>"01000", 469=>"01000", 
470=>"01000", 471=>"01000", 472=>"01000", 473=>"01000", 474=>"00101", 
475=>"00101", 476=>"00101", 477=>"00101", 478=>"00101", 479=>"00101", 
480=>"00101", 481=>"01000", 482=>"00101", 483=>"00101", 484=>"00101", 
485=>"00101", 486=>"01000", 487=>"01000", 488=>"01000", 489=>"00101", 
490=>"00101", 491=>"00101", 492=>"00101", 493=>"00101", 494=>"00101", 
495=>"00101", 496=>"00101", 497=>"00101", 498=>"00101", 499=>"00101", 
500=>"00101", 501=>"01000", 502=>"01000", 503=>"01000", 504=>"00101", 
505=>"00101", 506=>"00101", 507=>"00101", 508=>"00101", 509=>"00101", 
510=>"00101", 511=>"00101", 512=>"00101", 513=>"00101", 514=>"00101", 
515=>"00101", 516=>"00101", 517=>"00101", 518=>"00101", 519=>"00101", 
520=>"00101", 521=>"00101", 522=>"00101", 523=>"00101", 524=>"00101", 
525=>"00101", 526=>"00101", 527=>"00101", 528=>"00101", 529=>"00101", 
530=>"00101", 531=>"00101", 532=>"00101", 533=>"00101", 534=>"00101", 
535=>"00101", 536=>"00101", 537=>"00101", 538=>"00101", 539=>"00101", 
540=>"00101", 541=>"00101", 542=>"00101", 543=>"00101", 544=>"00101", 
545=>"00101", 546=>"00101", 547=>"00101", 548=>"00101", 549=>"00101", 
550=>"00101", 551=>"00101", 552=>"00101", 553=>"00101", 554=>"00101", 
555=>"00101", 556=>"00101", 557=>"00101", 558=>"00101", 559=>"00101", 
560=>"00101", 561=>"00101", 562=>"00101", 563=>"00101", 564=>"00101", 
565=>"00101", 566=>"00101", 567=>"00101", 568=>"00101", 569=>"00101", 
570=>"00101", 571=>"00101", 572=>"00101", 573=>"00101", 574=>"00101", 
575=>"00101", 576=>"00101", 577=>"00101", 578=>"00101", 579=>"00101", 
580=>"00101", 581=>"00101", 582=>"00101", 583=>"00101", 584=>"00101", 
585=>"00101", 586=>"00101", 587=>"00101", 588=>"00101", 589=>"00101", 
590=>"00101", 591=>"00101", 592=>"00101", 593=>"00101", 594=>"00101", 
595=>"00101", 596=>"00101", 597=>"00101", 598=>"00101", 599=>"00101", 
600=>"00101", 601=>"00101", 602=>"00101", 603=>"00101", 604=>"00101", 
605=>"00101", 606=>"00101", 607=>"00101", 608=>"00101", 609=>"00101", 
610=>"00101", 611=>"00101", 612=>"00101", 613=>"00101", 614=>"00101", 
615=>"00101", 616=>"00101", 617=>"00101", 618=>"00101", 619=>"00101", 
620=>"00101", 621=>"00101", 622=>"00101", 623=>"00101", 624=>"00101", 
625=>"00101", 626=>"00101", 627=>"00101", 628=>"00101", 629=>"00101", 
630=>"00101", 631=>"00101", 632=>"00101", 633=>"00101", 634=>"00101", 
635=>"00010", 636=>"00010", 637=>"00010", 638=>"00010", 639=>"00010", 
640=>"00010", 641=>"00010", 642=>"00101", 643=>"00101", 644=>"00101", 
645=>"00101", 646=>"00101", 647=>"00101", 648=>"00010", 649=>"00010", 
650=>"00010", 651=>"00010", 652=>"00010", 653=>"00010", 654=>"00010", 
655=>"00010", 656=>"00010", 657=>"00010", 658=>"00010", 659=>"00101", 
660=>"00101", 661=>"00101", 662=>"00010", 663=>"00010", 664=>"00010", 
665=>"00010", 666=>"00010", 667=>"00010", 668=>"00010", 669=>"00010", 
670=>"00010", 671=>"00010", 672=>"00010", 673=>"00010", 674=>"00010", 
675=>"00101", 676=>"00010", 677=>"00010", 678=>"00010", 679=>"00010", 
680=>"00010", 681=>"00010", 682=>"00010", 683=>"00010", 684=>"00010", 
685=>"00010", 686=>"00010", 687=>"00010", 688=>"00010", 689=>"00010", 
690=>"00010", 691=>"00010", 692=>"00010", 693=>"00010", 694=>"00010", 
695=>"00010", 696=>"00010", 697=>"00010", 698=>"00100", 699=>"00100", 
700=>"00010", 701=>"00010", 702=>"00010", 703=>"00010", 704=>"00010", 
705=>"00010", 706=>"00010", 707=>"00010", 708=>"00010", 709=>"00010", 
710=>"00010", 711=>"00010", 712=>"00010", 713=>"00010", 714=>"00010", 
715=>"00100", 716=>"00010", 717=>"00010", 718=>"00010", 719=>"00010", 
720=>"00010", 721=>"00010", 722=>"00010", 723=>"00010", 724=>"00100", 
725=>"00010", 726=>"00010", 727=>"00010", 728=>"00010", 729=>"00010", 
730=>"00100", 731=>"00100", 732=>"00100", 733=>"00010", 734=>"00010", 
735=>"00010", 736=>"00010", 737=>"00010", 738=>"00010", 739=>"00010", 
740=>"00010", 741=>"00010", 742=>"00010", 743=>"00010", 744=>"00010", 
745=>"00010", 746=>"00010", 747=>"00100", 748=>"00010", 749=>"00010", 
750=>"00010", 751=>"00010", 752=>"00010", 753=>"00010", 754=>"00010", 
755=>"00010", 756=>"00010", 757=>"00010", 758=>"00010", 759=>"00010", 
760=>"00010", 761=>"00010", 762=>"00100", 763=>"00010", 764=>"00010", 
765=>"00010", 766=>"00010", 767=>"00010", 768=>"00010", 769=>"00010", 
770=>"00010", 771=>"00010", 772=>"00010", 773=>"00010", 774=>"00010", 
775=>"00010", 776=>"00010", 777=>"00100", 778=>"00010", 779=>"00010", 
780=>"00010", 781=>"00010", 782=>"00010", 783=>"00010", 784=>"00010", 
785=>"00010", 786=>"00010", 787=>"00010", 788=>"00010", 789=>"00010", 
790=>"00010", 791=>"00010", 792=>"00100", 793=>"00010", 794=>"00010", 
795=>"00010", 796=>"00010", 797=>"00010", 798=>"00010", 799=>"00010", 
800=>"00010", 801=>"00010", 802=>"00010", 803=>"00010", 804=>"00010", 
805=>"00010", 806=>"00100", 807=>"00100", 808=>"00010", 809=>"00010", 
810=>"00010", 811=>"00010", 812=>"00010", 813=>"00010", 814=>"00100", 
815=>"00010", 816=>"00010", 817=>"00010", 818=>"00010", 819=>"00010", 
820=>"00100", 821=>"00100", 822=>"00010", 823=>"00010", 824=>"00010", 
825=>"00010", 826=>"00010", 827=>"00010", 828=>"00010", 829=>"00010", 
830=>"00010", 831=>"00010", 832=>"00010", 833=>"00010", 834=>"00010", 
835=>"00100", 836=>"00010", 837=>"00010", 838=>"00010", 839=>"00010", 
840=>"00010", 841=>"00010", 842=>"00010", 843=>"00010", 844=>"00010", 
845=>"00010", 846=>"00010", 847=>"00010", 848=>"00010", 849=>"00100", 
850=>"00100", 851=>"00010", 852=>"00010", 853=>"00010", 854=>"00010", 
855=>"00011", 856=>"00010", 857=>"00010", 858=>"00010", 859=>"00010", 
860=>"00010", 861=>"00010", 862=>"00010", 863=>"00010", 864=>"00100", 
865=>"00010", 866=>"00010", 867=>"00010", 868=>"00010", 869=>"00010", 
870=>"00011", 871=>"00011", 872=>"00010", 873=>"00010", 874=>"00010", 
875=>"00010", 876=>"00010", 877=>"00010", 878=>"00010", 879=>"00010", 
880=>"00010", 881=>"00010", 882=>"00010", 883=>"00010", 884=>"00010", 
885=>"00011", 886=>"00011", 887=>"00011", 888=>"00010", 889=>"00010", 
890=>"00010", 891=>"00010", 892=>"00010", 893=>"00010", 894=>"00010", 
895=>"00010", 896=>"00010", 897=>"00010", 898=>"00010", 899=>"00011", 
900=>"00011", 901=>"00011", 902=>"00011", 903=>"00011", 904=>"00011", 
905=>"00010", 906=>"00010", 907=>"00010", 908=>"00010", 909=>"00010", 
910=>"00010", 911=>"00010", 912=>"00011", 913=>"00011", 914=>"00011", 
915=>"00011", 916=>"00011", 917=>"00011", 918=>"00011", 919=>"00011", 
920=>"00011", 921=>"00011", 922=>"00011", 923=>"00011", 924=>"00011", 
925=>"00011", 926=>"00011", 927=>"00011", 928=>"00011", 929=>"00011", 
930=>"00011", 931=>"00011", 932=>"00011", 933=>"00011", 934=>"00011", 
935=>"00011", 936=>"00011", 937=>"00011", 938=>"00011", 939=>"00011", 
940=>"00011", 941=>"00011", 942=>"00011", 943=>"00011", 944=>"00011", 
945=>"00011", 946=>"00011", 947=>"00011", 948=>"00011", 949=>"00011", 
950=>"00011", 951=>"00011", 952=>"00011", 953=>"00011", 954=>"00011", 
955=>"00011", 956=>"00011", 957=>"00011", 958=>"00011", 959=>"00011", 
960=>"00011", 961=>"00011", 962=>"00011", 963=>"00011", 964=>"00011", 
965=>"00011", 966=>"00011", 967=>"00011", 968=>"00011", 969=>"00011", 
970=>"00011", 971=>"00011", 972=>"00011", 973=>"00011", 974=>"00011", 
975=>"00011", 976=>"00011", 977=>"00011", 978=>"00011", 979=>"00011", 
980=>"00011", 981=>"00011", 982=>"00011", 983=>"00011", 984=>"00011", 
985=>"00011", 986=>"00011", 987=>"00011", 988=>"00011", 989=>"00011", 
990=>"00011", 991=>"00011", 992=>"00011", 993=>"00011", 994=>"00011", 
995=>"00110", 996=>"00011", 997=>"00011", 998=>"00011", 999=>"00011", 
1000=>"00011", 1001=>"00011", 1002=>"00011", 1003=>"00011", 1004=>"00011", 
1005=>"00011", 1006=>"00011", 1007=>"00011", 1008=>"00011", 1009=>"00011", 
1010=>"00110", 1011=>"00110", 1012=>"00011", 1013=>"00011", 1014=>"00011", 
1015=>"00011", 1016=>"00011", 1017=>"00011", 1018=>"00011", 1019=>"00011", 
1020=>"00011", 1021=>"00011", 1022=>"00011", 1023=>"00011", 1024=>"00011", 
1025=>"00011", 1026=>"00110", 1027=>"00011", 1028=>"00011", 1029=>"00011", 
1030=>"00011", 1031=>"00011", 1032=>"00011", 1033=>"00011", 1034=>"00011", 
1035=>"00011", 1036=>"00011", 1037=>"00011", 1038=>"00011", 1039=>"00011", 
1040=>"00011", 1041=>"00110", 1042=>"00011", 1043=>"00011", 1044=>"00011", 
1045=>"00011", 1046=>"00011", 1047=>"00011", 1048=>"00011", 1049=>"00011", 
1050=>"00011", 1051=>"00011", 1052=>"00011", 1053=>"00011", 1054=>"00011", 
1055=>"00110", 1056=>"00110", 1057=>"00011", 1058=>"00011", 1059=>"00011", 
1060=>"00011", 1061=>"00011", 1062=>"00011", 1063=>"00011", 1064=>"00011", 
1065=>"00011", 1066=>"00011", 1067=>"00011", 1068=>"00011", 1069=>"00011", 
1070=>"00110", 1071=>"01000", 1072=>"00110", 1073=>"00110", 1074=>"00110", 
1075=>"00110", 1076=>"00110", 1077=>"00011", 1078=>"00011", 1079=>"00011", 
1080=>"00011", 1081=>"00011", 1082=>"00011", 1083=>"00011", 1084=>"00011", 
1085=>"00110", 1086=>"01000", 1087=>"01000", 1088=>"01000", 1089=>"01000", 
1090=>"01000", 1091=>"00110", 1092=>"00110", 1093=>"00011", 1094=>"00011", 
1095=>"00011", 1096=>"00011", 1097=>"00011", 1098=>"00011", 1099=>"00011", 
1100=>"00110", 1101=>"01000", 1102=>"01000", 1103=>"01000", 1104=>"01000", 
1105=>"01000", 1106=>"01000", 1107=>"00110", 1108=>"00011", 1109=>"00011", 
1110=>"00000", 1111=>"00000", 1112=>"00000", 1113=>"00000", 1114=>"00000", 
1115=>"00110", 1116=>"01000", 1117=>"01000", 1118=>"01000", 1119=>"01000", 
1120=>"01000", 1121=>"01000", 1122=>"01000", 1123=>"00000", 1124=>"00000", 
1125=>"01000", 1126=>"01000", 1127=>"01000", 1128=>"01000", 1129=>"01000", 
1130=>"00110", 1131=>"01000", 1132=>"01000", 1133=>"01000", 1134=>"01000", 
1135=>"01000", 1136=>"01000", 1137=>"01000", 1138=>"01000", 1139=>"01000", 
1140=>"01000", 1141=>"01000", 1142=>"01000", 1143=>"01000", 1144=>"01000", 
1145=>"01000", 1146=>"01000", 1147=>"01000", 1148=>"01000", 1149=>"01000", 
1150=>"01000", 1151=>"01000", 1152=>"01000", 1153=>"01000", 1154=>"01000", 
1155=>"01000", 1156=>"01000", 1157=>"01000", 1158=>"01000", 1159=>"01000", 
1160=>"01000", 1161=>"01000", 1162=>"01000", 1163=>"01000", 1164=>"01000", 
1165=>"01000", 1166=>"01000", 1167=>"01000", 1168=>"01000", 1169=>"01000", 
1170=>"01000", 1171=>"01000", 1172=>"01000", 1173=>"01000", 1174=>"01000", 
1175=>"01000", 1176=>"01000", 1177=>"01000", 1178=>"01000", 1179=>"01000", 
1180=>"01000", 1181=>"01000", 1182=>"01000", 1183=>"01000", 1184=>"01000", 
1185=>"01000", 1186=>"01000", 1187=>"01000", 1188=>"01000", 1189=>"01000", 
1190=>"01000", 1191=>"01000", 1192=>"01000", 1193=>"00110", 1194=>"00110", 
1195=>"00110", 1196=>"01000", 1197=>"01000", 1198=>"01000", 1199=>"01000", 
1200=>"01000", 1201=>"01000", 1202=>"01000", 1203=>"01000", 1204=>"01000", 
1205=>"01000", 1206=>"01000", 1207=>"00110", 1208=>"00110", 1209=>"00111", 
1210=>"00110", 1211=>"01000", 1212=>"01000", 1213=>"01000", 1214=>"01000", 
1215=>"01000", 1216=>"01000", 1217=>"01000", 1218=>"01000", 1219=>"01000", 
1220=>"00110", 1221=>"00110", 1222=>"00111", 1223=>"00111", 1224=>"00111", 
1225=>"00110", 1226=>"00110", 1227=>"00110", 1228=>"01000", 1229=>"01000", 
1230=>"01000", 1231=>"01000", 1232=>"01000", 1233=>"01000", 1234=>"01000", 
1235=>"01000", 1236=>"00110", 1237=>"00111", 1238=>"00111", 1239=>"00111", 
1240=>"00111", 1241=>"00111", 1242=>"00110", 1243=>"01000", 1244=>"01000", 
1245=>"01000", 1246=>"01000", 1247=>"01000", 1248=>"01000", 1249=>"01000", 
1250=>"01000", 1251=>"00110", 1252=>"00111", 1253=>"00111", 1254=>"00111", 
1255=>"00111", 1256=>"00110", 1257=>"00110", 1258=>"01000", 1259=>"01000", 
1260=>"01000", 1261=>"01000", 1262=>"01000", 1263=>"01000", 1264=>"01000", 
1265=>"01000", 1266=>"00110", 1267=>"00110", 1268=>"00110", 1269=>"00110", 
1270=>"00110", 1271=>"00110", 1272=>"01000", 1273=>"01000", 1274=>"01000", 
1275=>"01000", 1276=>"01000", 1277=>"01000", 1278=>"01000", 1279=>"01000", 
1280=>"01000", 1281=>"01000", 1282=>"01000", 1283=>"01000", 1284=>"01000", 
1285=>"01000", 1286=>"01000", 1287=>"01000", 1288=>"01000", 1289=>"01000", 
1290=>"01000", 1291=>"01000", 1292=>"01000", 1293=>"01000", 1294=>"01000", 
1295=>"01000", 1296=>"01000", 1297=>"01000", 1298=>"01000", 1299=>"01000", 
1300=>"01000", 1301=>"01000", 1302=>"01000", 1303=>"01000", 1304=>"01000", 
1305=>"01000", 1306=>"01000", 1307=>"01000", 1308=>"01000", 1309=>"01000", 
1310=>"01000", 1311=>"01000", 1312=>"00110", 1313=>"00110", 1314=>"00110", 
1315=>"00110", 1316=>"00110", 1317=>"00110", 1318=>"01000", 1319=>"01000", 
1320=>"01000", 1321=>"01000", 1322=>"01000", 1323=>"01000", 1324=>"01000", 
1325=>"01000", 1326=>"01000", 1327=>"00110", 1328=>"00110", 1329=>"01000", 
1330=>"01000", 1331=>"01000", 1332=>"01000", 1333=>"01000", 1334=>"01000", 
1335=>"01000", 1336=>"01000", 1337=>"01000", 1338=>"01000", 1339=>"01000", 
1340=>"01000", 1341=>"01000", 1342=>"01000", 1343=>"00110", 1344=>"00110", 
1345=>"00110", 1346=>"01000", 1347=>"01000", 1348=>"01000", 1349=>"01000", 
1350=>"01000", 1351=>"01000", 1352=>"01000", 1353=>"01000", 1354=>"01000", 
1355=>"01000", 1356=>"01000", 1357=>"01000", 1358=>"01000", 1359=>"01000", 
1360=>"00110", 1361=>"00110", 1362=>"01000", 1363=>"01000", 1364=>"01000", 
1365=>"01000", 1366=>"01000", 1367=>"01000", 1368=>"01000", 1369=>"01000", 
1370=>"01000", 1371=>"01000", 1372=>"01000", 1373=>"01000", 1374=>"01000", 
1375=>"01000", 1376=>"00110", 1377=>"01000", 1378=>"01000", 1379=>"01000", 
1380=>"01000", 1381=>"01000", 1382=>"01000", 1383=>"01000", 1384=>"01000", 
1385=>"01000", 1386=>"01000", 1387=>"01000", 1388=>"01000", 1389=>"01000", 
1390=>"01000", 1391=>"00110", 1392=>"01000", 1393=>"01000", 1394=>"01000", 
1395=>"01000", 1396=>"01000", 1397=>"01000", 1398=>"01000", 1399=>"01000", 
1400=>"01000", 1401=>"01000", 1402=>"00110", 1403=>"00110", 1404=>"00110", 
1405=>"00110", 1406=>"00110", 1407=>"01000", 1408=>"01000", 1409=>"01000", 
1410=>"01000", 1411=>"01000", 1412=>"01000", 1413=>"01000", 1414=>"01000", 
1415=>"01000", 1416=>"01000", 1417=>"00110", 1418=>"01000", 1419=>"01000", 
1420=>"01000", 1421=>"01000", 1422=>"01000", 1423=>"01000", 1424=>"01000", 
1425=>"01000", 1426=>"01000", 1427=>"01000", 1428=>"01000", 1429=>"01000", 
1430=>"01000", 1431=>"01000", 1432=>"01000", 1433=>"01000", 1434=>"01000", 
1435=>"01000", 1436=>"01000", 1437=>"01000", 1438=>"01000", 1439=>"01000", 
1440=>"01000", 1441=>"01000", 1442=>"01000", 1443=>"00001", 1444=>"00001", 
1445=>"00001", 1446=>"00001", 1447=>"00001", 1448=>"01000", 1449=>"01000", 
1450=>"01000", 1451=>"01000", 1452=>"01000", 1453=>"01000", 1454=>"01000", 
1455=>"01000", 1456=>"00001", 1457=>"00001", 1458=>"00001", 1459=>"00001", 
1460=>"00001", 1461=>"00001", 1462=>"00001", 1463=>"00001", 1464=>"00001", 
1465=>"00001", 1466=>"01000", 1467=>"01000", 1468=>"01000", 1469=>"01000", 
1470=>"00001", 1471=>"00001", 1472=>"00001", 1473=>"00001", 1474=>"00001", 
1475=>"00001", 1476=>"00001", 1477=>"00001", 1478=>"00001", 1479=>"00001", 
1480=>"00001", 1481=>"00001", 1482=>"00001", 1483=>"01000", 1484=>"01000", 
1485=>"00001", 1486=>"00001", 1487=>"00001", 1488=>"00001", 1489=>"00001", 
1490=>"00001", 1491=>"00001", 1492=>"00001", 1493=>"00001", 1494=>"00001", 
1495=>"00001", 1496=>"00001", 1497=>"00001", 1498=>"01000", 1499=>"01000", 
1500=>"00001", 1501=>"00001", 1502=>"00001", 1503=>"00001", 1504=>"00001", 
1505=>"00001", 1506=>"00001", 1507=>"00001", 1508=>"00001", 1509=>"00001", 
1510=>"00001", 1511=>"00001", 1512=>"00001", 1513=>"00001", 1514=>"01000", 
1515=>"00001", 1516=>"00001", 1517=>"00001", 1518=>"00001", 1519=>"00001", 
1520=>"00001", 1521=>"00001", 1522=>"00001", 1523=>"00001", 1524=>"01000", 
1525=>"01000", 1526=>"01000", 1527=>"01000", 1528=>"00001", 1529=>"01000", 
1530=>"00001", 1531=>"00001", 1532=>"00001", 1533=>"00001", 1534=>"00001", 
1535=>"00001", 1536=>"00001", 1537=>"01000", 1538=>"01000", 1539=>"01000", 
1540=>"01000", 1541=>"00001", 1542=>"00001", 1543=>"00001", 1544=>"01000", 
1545=>"00001", 1546=>"00001", 1547=>"00001", 1548=>"00001", 1549=>"00001", 
1550=>"00001", 1551=>"01000", 1552=>"01000", 1553=>"01000", 1554=>"01000", 
1555=>"01000", 1556=>"00001", 1557=>"00001", 1558=>"00001", 1559=>"01000", 
1560=>"00001", 1561=>"00001", 1562=>"00001", 1563=>"00001", 1564=>"00001", 
1565=>"00001", 1566=>"01000", 1567=>"01000", 1568=>"01000", 1569=>"01000", 
1570=>"01000", 1571=>"00001", 1572=>"00001", 1573=>"00001", 1574=>"01000", 
1575=>"00001", 1576=>"00001", 1577=>"00001", 1578=>"00001", 1579=>"00001", 
1580=>"00001", 1581=>"00001", 1582=>"00001", 1583=>"01000", 1584=>"01000", 
1585=>"01000", 1586=>"00001", 1587=>"00001", 1588=>"00001", 1589=>"01000", 
1590=>"00001", 1591=>"00001", 1592=>"00001", 1593=>"00001", 1594=>"00001", 
1595=>"00001", 1596=>"00001", 1597=>"00001", 1598=>"00001", 1599=>"00001", 
1600=>"01000", 1601=>"01000", 1602=>"00001", 1603=>"00001", 1604=>"01000", 
1605=>"00001", 1606=>"00001", 1607=>"00001", 1608=>"00001", 1609=>"00001", 
1610=>"00001", 1611=>"00001", 1612=>"00001", 1613=>"00001", 1614=>"00001", 
1615=>"00001", 1616=>"01000", 1617=>"01000", 1618=>"01000", 1619=>"01000", 
1620=>"01000", 1621=>"00001", 1622=>"00001", 1623=>"00001", 1624=>"00001", 
1625=>"00001", 1626=>"00001", 1627=>"00001", 1628=>"00001", 1629=>"00001", 
1630=>"00001", 1631=>"00001", 1632=>"01000", 1633=>"00110", 1634=>"01000", 
1635=>"01000", 1636=>"01000", 1637=>"00001", 1638=>"00001", 1639=>"00001", 
1640=>"00001", 1641=>"00001", 1642=>"00001", 1643=>"00001", 1644=>"00001", 
1645=>"00001", 1646=>"01000", 1647=>"01000", 1648=>"01000", 1649=>"01000", 
1650=>"01000", 1651=>"01000", 1652=>"01000", 1653=>"00001", 1654=>"00001", 
1655=>"00001", 1656=>"00001", 1657=>"01000", 1658=>"00001", 1659=>"00001", 
1660=>"01000", 1661=>"01000", 1662=>"01000", 1663=>"01000", 1664=>"01000", 
1665=>"01000", 1666=>"01000", 1667=>"01000", 1668=>"01000", 1669=>"01000", 
1670=>"01000", 1671=>"01000", 1672=>"01000", 1673=>"01000", 1674=>"01000", 
1675=>"01000", 1676=>"01000", 1677=>"01000", 1678=>"01000", 1679=>"01000", 
1680=>"01000", 1681=>"01000", 1682=>"01000", 1683=>"01000", 1684=>"01000", 
1685=>"01000", 1686=>"01000", 1687=>"00110", 1688=>"01000", 1689=>"01000", 
1690=>"01000", 1691=>"01000", 1692=>"01000", 1693=>"01000", 1694=>"01000", 
1695=>"01000", 1696=>"01000", 1697=>"01000", 1698=>"01000", 1699=>"01000", 
1700=>"01000", 1701=>"01000", 1702=>"00110", 1703=>"01000", 1704=>"01000", 
1705=>"01000", 1706=>"01000", 1707=>"01000", 1708=>"01000", 1709=>"01000", 
1710=>"01000", 1711=>"01000", 1712=>"01000", 1713=>"01000", 1714=>"01000", 
1715=>"01000", 1716=>"00110", 1717=>"00110", 1718=>"00110", 1719=>"00110", 
1720=>"00110", 1721=>"00110", 1722=>"00110", 1723=>"00110", 1724=>"01000", 
1725=>"01000", 1726=>"01000", 1727=>"01000", 1728=>"01000", 1729=>"01000", 
1730=>"01000", 1731=>"01000", 1732=>"00110", 1733=>"01000", 1734=>"01000", 
1735=>"01000", 1736=>"01000", 1737=>"01000", 1738=>"01000", 1739=>"01000", 
1740=>"01000", 1741=>"01000", 1742=>"01000", 1743=>"01000", 1744=>"01000", 
1745=>"01000", 1746=>"01000", 1747=>"00110", 1748=>"01000", 1749=>"01000", 
1750=>"01000", 1751=>"01000", 1752=>"01000", 1753=>"01000", 1754=>"01000", 
1755=>"01000", 1756=>"01000", 1757=>"01000", 1758=>"01000", 1759=>"01000", 
1760=>"01000", 1761=>"01000", 1762=>"00110", 1763=>"01000", 1764=>"01000", 
1765=>"01000", 1766=>"01000", 1767=>"01000", 1768=>"01000", 1769=>"01000", 
1770=>"01000", 1771=>"01000", 1772=>"01000", 1773=>"01000", 1774=>"01000", 
1775=>"01000", 1776=>"01000", 1777=>"01000", 1778=>"01000", 1779=>"01000", 
1780=>"01000", 1781=>"01000", 1782=>"01000", 1783=>"01000", 1784=>"01000", 
1785=>"01000", 1786=>"01000", 1787=>"01000", 1788=>"01000", 1789=>"01000", 
1790=>"01000", 1791=>"01000", 1792=>"01000", 1793=>"01000", 1794=>"01000", 
1795=>"01000", 1796=>"01000", 1797=>"01000", 1798=>"01000", 1799=>"01000", 
1800=>"01000", 1801=>"01000", 1802=>"01000", 1803=>"01000", 1804=>"01000", 
1805=>"01000", 1806=>"01000", 1807=>"01000", 1808=>"01000", 1809=>"01000", 
1810=>"01000", 1811=>"01000", 1812=>"01000", 1813=>"01000", 1814=>"01000", 
1815=>"01000", 1816=>"01000", 1817=>"01000", 1818=>"01000", 1819=>"01000", 
1820=>"01000", 1821=>"01000", 1822=>"01000", 1823=>"01000", 1824=>"01000", 
1825=>"01000", 1826=>"01000", 1827=>"01000", 1828=>"01000", 1829=>"01000", 
1830=>"01000", 1831=>"01000", 1832=>"01000", 1833=>"01000", 1834=>"01000", 
1835=>"01000", 1836=>"01000", 1837=>"01000", 1838=>"01000", 1839=>"01000", 
1840=>"01000", 1841=>"01000", 1842=>"01000", 1843=>"01000", 1844=>"01000", 
1845=>"01000", 1846=>"01000", 1847=>"01000", 1848=>"01000", 1849=>"01000", 
1850=>"01000", 1851=>"01000", 1852=>"01000", 1853=>"01000", 1854=>"01000", 
1855=>"01000", 1856=>"01000", 1857=>"01000", 1858=>"01000", 1859=>"01000", 
1860=>"01000", 1861=>"01000", 1862=>"01000", 1863=>"01000", 1864=>"01000", 
1865=>"01000", 1866=>"01000", 1867=>"01000", 1868=>"01000", 1869=>"01000", 
1870=>"01000", 1871=>"01000", 1872=>"01000", 1873=>"01000", 1874=>"01000", 
1875=>"01000", 1876=>"01000", 1877=>"01000", 1878=>"01000", 1879=>"01000", 
1880=>"01000", 1881=>"01000", 1882=>"01000", 1883=>"01000", 1884=>"01000", 
1885=>"01000", 1886=>"01000", 1887=>"01000", 1888=>"01000", 1889=>"01000", 
1890=>"01000", 1891=>"01000", 1892=>"01000", 1893=>"01000", 1894=>"01000", 
1895=>"01000", 1896=>"01000", 1897=>"01000", 1898=>"01000", 1899=>"01000", 
1900=>"01000", 1901=>"01000", 1902=>"01000", 1903=>"01000", 1904=>"01000", 
1905=>"01000", 1906=>"01000", 1907=>"01000", 1908=>"01000", 1909=>"01000", 
1910=>"01000", 1911=>"01000", 1912=>"01000", 1913=>"01000", 1914=>"01000", 
1915=>"01000", 1916=>"01000", 1917=>"01000", 1918=>"01000", 1919=>"01000", 
1920=>"01000", 1921=>"01000", 1922=>"01000", 1923=>"01000", 1924=>"01000", 
1925=>"01000", 1926=>"01000", 1927=>"01000", 1928=>"01000", 1929=>"01000", 
1930=>"01000", 1931=>"01000", 1932=>"01000", 1933=>"01000", 1934=>"01000", 
1935=>"01000", 1936=>"01000", 1937=>"01000", 1938=>"01000", 1939=>"01000", 
1940=>"01000", 1941=>"01000", 1942=>"01000", 1943=>"01000", 1944=>"01000", 
1945=>"01000", 1946=>"01000", 1947=>"01000", 1948=>"01000", 1949=>"01000", 
1950=>"01000", 1951=>"01000", 1952=>"01000", 1953=>"01000", 1954=>"01000", 
1955=>"01000", 1956=>"01000", 1957=>"01000", 1958=>"01000", 1959=>"01000", 
1960=>"01000", 1961=>"01000", 1962=>"01000", 1963=>"01000", 1964=>"01000", 
1965=>"01000", 1966=>"01000", 1967=>"01000", 1968=>"01000", 1969=>"01000", 
1970=>"01000", 1971=>"01000", 1972=>"01000", 1973=>"01000", 1974=>"01000", 
1975=>"01000", 1976=>"01000", 1977=>"01000", 1978=>"01000", 1979=>"01000", 
1980=>"01000", 1981=>"01000", 1982=>"01000", 1983=>"01000", 1984=>"01000", 
1985=>"01000", 1986=>"01000", 1987=>"01000", 1988=>"01000", 1989=>"01000", 
1990=>"01000", 1991=>"01000", 1992=>"01000", 1993=>"01000", 1994=>"01000", 
1995=>"01000", 1996=>"01000", 1997=>"01000", 1998=>"01000", 1999=>"01000", 
2000=>"01000", 2001=>"01000", 2002=>"01000", 2003=>"01000", 2004=>"01000", 
2005=>"01000", 2006=>"01000", 2007=>"01000", 2008=>"01000", 2009=>"01000", 
2010=>"01000", 2011=>"01000", 2012=>"01000", 2013=>"01000", 2014=>"01000", 
2015=>"01000", 2016=>"01000", 2017=>"01000", 2018=>"01000", 2019=>"01000", 
2020=>"01000", 2021=>"01000", 2022=>"01000", 2023=>"01000", 2024=>"01000", 
2025=>"01000", 2026=>"01000", 2027=>"01000", 2028=>"01000", 2029=>"01000", 
2030=>"01000", 2031=>"01000", 2032=>"01000", 2033=>"01000", 2034=>"01000", 
2035=>"01000", 2036=>"01000", 2037=>"01000", 2038=>"01000", 2039=>"01000", 
2040=>"01000", 2041=>"01000", 2042=>"01000", 2043=>"01000", 2044=>"01000", 
2045=>"01000", 2046=>"01000", 2047=>"01000", 2048=>"01000", 2049=>"01000", 
2050=>"01000", 2051=>"01000", 2052=>"01000", 2053=>"01000", 2054=>"01000", 
2055=>"01000", 2056=>"01000", 2057=>"01000", 2058=>"01000", 2059=>"01000", 
2060=>"01000", 2061=>"01000", 2062=>"01000", 2063=>"01000", 2064=>"01000", 
2065=>"01000", 2066=>"01000", 2067=>"01000", 2068=>"01000", 2069=>"01000", 
2070=>"01000", 2071=>"01000", 2072=>"01000", 2073=>"01000", 2074=>"01000", 
2075=>"01000", 2076=>"01000", 2077=>"01000", 2078=>"01000", 2079=>"01000", 
2080=>"01000", 2081=>"01000", 2082=>"01000", 2083=>"01000", 2084=>"01000", 
2085=>"01000", 2086=>"01000", 2087=>"01000", 2088=>"01000", 2089=>"01000", 
2090=>"01000", 2091=>"01000", 2092=>"01000", 2093=>"01000", 2094=>"01000", 
2095=>"01000", 2096=>"01000", 2097=>"01000", 2098=>"01000", 2099=>"01000", 
2100=>"01000", 2101=>"01000", 2102=>"01000", 2103=>"01000", 2104=>"01000", 
2105=>"01000", 2106=>"01000", 2107=>"01000", 2108=>"01000", 2109=>"01000", 
2110=>"01000", 2111=>"01000", 2112=>"01000", 2113=>"01000", 2114=>"01000", 
2115=>"01000", 2116=>"01000", 2117=>"01000", 2118=>"01000", 2119=>"01000", 
2120=>"01000", 2121=>"01000", 2122=>"01000", 2123=>"01000", 2124=>"01000", 
2125=>"01000", 2126=>"01000", 2127=>"01000", 2128=>"01000", 2129=>"01000", 
2130=>"01000", 2131=>"01000", 2132=>"01000", 2133=>"01000", 2134=>"01000", 
2135=>"01000", 2136=>"01000", 2137=>"01000", 2138=>"01000", 2139=>"01000", 
2140=>"01000", 2141=>"01000", 2142=>"01000", 2143=>"01000", 2144=>"01000", 
2145=>"01000", 2146=>"01000", 2147=>"01000", 2148=>"01000", 2149=>"01000", 
2150=>"01000", 2151=>"01000", 2152=>"01000", 2153=>"01000", 2154=>"01000", 
2155=>"01000", 2156=>"01000", 2157=>"01000", 2158=>"01000", 2159=>"01000", 
2160=>"01000", 2161=>"01000", 2162=>"01000", 2163=>"01000", 2164=>"01000", 
2165=>"01000", 2166=>"01000", 2167=>"01000", 2168=>"01000", 2169=>"01000", 
2170=>"01000", 2171=>"01000", 2172=>"01000", 2173=>"01000", 2174=>"01000", 
2175=>"01000", 2176=>"01000", 2177=>"01000", 2178=>"01000", 2179=>"01000", 
2180=>"01000", 2181=>"01000", 2182=>"01000", 2183=>"01000", 2184=>"01000", 
2185=>"01000", 2186=>"01000", 2187=>"01000", 2188=>"01000", 2189=>"01000", 
2190=>"01000", 2191=>"01000", 2192=>"01000", 2193=>"01000", 2194=>"01000", 
2195=>"01000", 2196=>"01000", 2197=>"01000", 2198=>"01000", 2199=>"01000", 
2200=>"01000", 2201=>"01000", 2202=>"01000", 2203=>"01000", 2204=>"01000", 
2205=>"01000", 2206=>"01000", 2207=>"01000", 2208=>"01000", 2209=>"01000", 
2210=>"01000", 2211=>"01000", 2212=>"01000", 2213=>"01000", 2214=>"01000", 
2215=>"01000", 2216=>"01000", 2217=>"01000", 2218=>"01000", 2219=>"01000", 
2220=>"01000", 2221=>"01000", 2222=>"01000", 2223=>"01000", 2224=>"01000", 
2225=>"01000", 2226=>"01000", 2227=>"01000", 2228=>"01000", 2229=>"01000", 
2230=>"01000", 2231=>"01000", 2232=>"01000", 2233=>"01000", 2234=>"01000", 
2235=>"01000", 2236=>"01000", 2237=>"01000", 2238=>"01000", 2239=>"01000", 
2240=>"01000", 2241=>"01000", 2242=>"01000", 2243=>"01000", 2244=>"01000", 
2245=>"01000", 2246=>"01000", 2247=>"01000", 2248=>"01000", 2249=>"01000" 

);

signal query_help : std_logic_vector(4 downto 0);

begin

    process(clk)
    begin
        if rising_edge(clk) then
            data_out <= pictMem(to_integer(addr));
			query_help <= pictMem(to_integer(query_addr));
        end if;
    end process;

	query_result <= '1' when query_help > 4 else '0';

end Behavioral;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity level_mem is
    port (
        clk      : in std_logic;
        data_out : out std_logic_vector(4 downto 0);
        addr    : in unsigned(11 downto 0);
		level_choice : in std_logic;
        query_addr : in unsigned(11 downto 0);
        query_result : out std_logic
         );
end level_mem;

architecture Behavioral of level_mem is
    type ram_t is array (0 to 2249) of std_logic_vector(4 downto 0);
    signal pictMem : ram_t := (
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "01010", "11111", "01000", "00000", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "01010", 
           "10010", "11111", "10101", "00111", "00000", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "01010", "10010", "11111", 
           "10010", "10010", "10010", "00100", "01001", 
           "11111", "11111", "11111", "11111", "11111", 
           "01010", "11111", "10010", "10110", "10010", 
           "10110", "10110", "10110", "00100", "00000", 
           "11111", "11111", "11111", "01010", "11111", 
           "11111", "10010", "10110", "10110", "10110", 
           "10110", "10110", "10110", "00100", "01001", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "10010", "10110", "10010", 
           "10110", "10110", "10110", "00100", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "10010", "11111", 
           "10010", "10010", "10010", "00100", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "10010", "11111", "11111", "00111", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "00111", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "00111", "01001", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "00111", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "00111", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "10101", "00111", "01001", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "00111", "01001", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "00010", "00000", "01001", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "00010", "00000", "01001", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "00010", "10101", "00111", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "00010", "10001", "00111", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "00010", "10000", "11111", "00111", "01001", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "00010", "11111", "11111", "00111", "01001", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "01000", 
           "01001", "01001", "01001", "00000", "01001", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "01000", 
           "11111", "11111", "11111", "00111", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "01000", "10000", "11111", "00111", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "01000", "11111", "11111", "00111", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "01000", "11111", "11111", "00111", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "01000", "10001", "11111", "00111", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "01000", "11111", "11111", "00111", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "01000", "11111", "11111", "00111", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "01000", 
           "11111", "11111", "11111", "00111", "01001", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "01000", 
           "01001", "11111", "11111", "00111", "01001", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "00010", "10001", "11111", "00111", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "00010", "10000", "11111", "00111", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "00010", "11111", "00111", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "00010", "10001", "00111", "01001", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "00010", "00111", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "00010", "00111", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "00111", "01001", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "00111", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "10101", "00111", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "00111", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "10101", "00111", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "00111", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "00111", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "00111", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "00011", "10000", "11111", 
           "11111", "11111", "10101", "00111", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "00011", "10010", "10010", "10010", 
           "10010", "10010", "10010", "00011", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "00011", "10110", "10110", "10110", "10110", 
           "10110", "10110", "10110", "00011", "00000", 
           "11111", "01010", "11111", "11111", "00011", 
           "10110", "10110", "10110", "10110", "10110", 
           "10110", "00100", "10110", "00011", "00000", 
           "11111", "01010", "11111", "00011", "10110", 
           "10110", "10110", "10110", "10110", "10110", 
           "10110", "00100", "10110", "00011", "00000", 
           "11111", "01010", "00011", "10110", "10110", 
           "10110", "10110", "10110", "10110", "10110", 
           "10110", "00100", "10110", "00011", "00000", 
           "11111", "00011", "10110", "10110", "10010", 
           "10010", "10010", "10010", "10110", "10110", 
           "10110", "00100", "10110", "00011", "00000", 
           "11111", "00011", "10110", "10110", "10010", 
           "11111", "11111", "10010", "10110", "10110", 
           "10110", "00100", "10110", "00011", "00000", 
           "11111", "00011", "10110", "10110", "10010", 
           "11111", "11111", "10010", "10110", "10110", 
           "10110", "10110", "10110", "00011", "00000", 
           "11111", "00011", "10110", "10110", "10010", 
           "10010", "10010", "10010", "10110", "10110", 
           "10110", "10110", "10110", "00011", "00000", 
           "11111", "00011", "10110", "10110", "10110", 
           "10110", "10110", "10110", "10110", "10110", 
           "00100", "10110", "10110", "00011", "00011", 
           "11111", "00011", "10110", "10110", "10110", 
           "10110", "10110", "10110", "10110", "10110", 
           "10110", "00100", "10110", "10110", "10110", 
           "11111", "00011", "10110", "10110", "10110", 
           "10110", "10110", "10110", "10110", "10110", 
           "10110", "00100", "10110", "10110", "10110", 
           "11111", "00011", "10110", "10110", "10110", 
           "10110", "10110", "10110", "10110", "10110", 
           "10110", "00100", "10110", "10110", "10110", 
           "11111", "00011", "10110", "10110", "10110", 
           "10110", "10110", "10110", "10110", "10110", 
           "10110", "00100", "10110", "10110", "10110", 
           "11111", "00011", "10110", "10110", "10110", 
           "10110", "10110", "10110", "10110", "10110", 
           "00100", "10110", "10110", "00011", "00011", 
           "11111", "00011", "10110", "10110", "10010", 
           "10010", "10010", "10010", "10110", "10110", 
           "10110", "10110", "10110", "00011", "00000", 
           "11111", "00011", "10110", "10110", "10010", 
           "11111", "11111", "10010", "10110", "10110", 
           "00100", "10110", "10110", "00011", "00000", 
           "11111", "00011", "10110", "10110", "10010", 
           "11111", "11111", "10010", "10110", "10110", 
           "00100", "10110", "00100", "00011", "00000", 
           "11111", "00011", "10110", "10110", "10010", 
           "10010", "10010", "10010", "10110", "10110", 
           "10110", "10110", "00100", "00011", "00000", 
           "11111", "00011", "10110", "10110", "10110", 
           "10110", "10110", "10110", "10110", "10110", 
           "10110", "10110", "10110", "00011", "00000", 
           "11111", "00011", "10110", "10110", "10110", 
           "10110", "10110", "10110", "10110", "00100", 
           "10110", "10110", "10110", "00011", "00000", 
           "11111", "00011", "10110", "10110", "10110", 
           "10110", "10110", "10110", "10110", "10110", 
           "10110", "10110", "10110", "00011", "00000", 
           "11111", "00011", "10110", "10110", "10110", 
           "10110", "10110", "10110", "10110", "10110", 
           "10110", "10110", "10110", "00011", "00000", 
           "11111", "00011", "10110", "10110", "10110", 
           "10110", "10110", "10110", "00100", "10110", 
           "10110", "10110", "10110", "00011", "00000", 
           "11111", "00011", "10110", "10110", "10110", 
           "10110", "10110", "10110", "10110", "10110", 
           "10110", "10110", "10110", "00011", "00000", 
           "11111", "00011", "10110", "10110", "10110", 
           "10110", "10110", "10110", "10110", "10110", 
           "10110", "10110", "10110", "00011", "00000", 
           "11111", "00011", "10110", "10110", "10110", 
           "10110", "10110", "10110", "00100", "10110", 
           "10110", "10110", "10110", "00011", "00000", 
           "11111", "00011", "10110", "10110", "10110", 
           "10110", "10110", "10110", "10110", "10110", 
           "10110", "10110", "10110", "00011", "00000", 
           "11111", "00011", "10110", "10110", "10110", 
           "10110", "10110", "10110", "10110", "10110", 
           "10110", "10110", "10110", "00011", "00000", 
           "11111", "00011", "10110", "10110", "10110", 
           "10110", "10110", "10110", "00100", "10110", 
           "10110", "10110", "10110", "00011", "00000", 
           "11111", "00011", "10110", "10110", "10110", 
           "10110", "10110", "10110", "10110", "10110", 
           "10110", "10110", "10110", "00011", "00000", 
           "11111", "01010", "00011", "10110", "10110", 
           "10110", "10110", "10110", "10110", "10110", 
           "10110", "10110", "10110", "00011", "00000", 
           "11111", "01010", "11111", "00011", "10110", 
           "10110", "10110", "00100", "10110", "10110", 
           "10110", "10110", "10110", "00011", "00000", 
           "11111", "01010", "11111", "11111", "10010", 
           "10110", "10110", "00100", "10110", "10110", 
           "10110", "10110", "10110", "00011", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "10010", "10110", "10110", "10110", "10110", 
           "10110", "10110", "10110", "00011", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "10010", "00100", "00100", "00100", 
           "00100", "00100", "00100", "00011", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "00100", "11111", "00011", "11111", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "00100", "00011", "11111", "11111", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "00100", "10000", "11111", "11111", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "00100", "11111", "11111", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "00100", "11111", "11111", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "00100", "11111", "11111", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "00100", "11111", "11111", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "00100", "11111", "11111", "11111", 
           "10011", "00001", "11111", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "00001", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "10011", "00001", "11111", "11111", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "00001", "11111", "11111", "11111", "11111", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "10011", "00001", "11111", "11111", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "10011", "00001", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "00001", "00000", "00000", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "10011", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "10011", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "00001", "00000", "00000", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "10011", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "01001", "01001", "00000", "00000", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "01001", "00000", "00000", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "01001", "00000", "00000", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "01001", "00000", "00000", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "01001", "00000", "00000", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "01001", "01001", "00000", "00000", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "00001", "00000", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "01001", "00000", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "00011", "00011", "00000", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "00011", "00011", "00011", "00000", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "00011", "00011", "00011", "00000", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "00011", "00000", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "00011", "00011", "00011", "00000", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "00011", "11111", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "00011", "11111", "11111", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "00011", 
           "10010", "10010", "10010", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "00011", "10010", 
           "10110", "10110", "10110", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "11111", "00011", "10010", "10110", 
           "10110", "10110", "10110", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "00011", "10010", "10110", "10110", 
           "10110", "10110", "10110", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "00011", "10010", "10110", "10110", 
           "10110", "10110", "10110", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "00011", "10010", "10110", "10110", 
           "10110", "10110", "10110", "00001", "00000", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "00011", "10010", "10110", "10110", 
           "10110", "10110", "10110", "00001", "00000", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "00011", "10010", "10010", "10010", 
           "10010", "10010", "10010", "00001", "00000");

signal you_win : ram_t := (
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "01010", "11111", "11111", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "01010", 
           "11111", "11111", "10011", "00001", "00000", 
           "11111", "11111", "11111", "11111", "11111", 
           "01010", "11111", "11111", "11111", "11111", 
           "11111", "01010", "11111", "00001", "00000", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "10010", "10010", "11111", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "10010", "11111", "11111", "11111", 
           "11111", "01010", "11111", "11111", "10010", 
           "10010", "11111", "10011", "00001", "00000", 
           "11111", "11111", "10010", "11111", "11111", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "10010", "11111", "00001", "00000", 
           "11111", "11111", "11111", "10010", "10010", 
           "10010", "01010", "11111", "11111", "11111", 
           "10010", "11111", "11111", "00001", "00000", 
           "11111", "11111", "10010", "11111", "11111", 
           "11111", "01010", "11111", "11111", "11111", 
           "11111", "10010", "11111", "00001", "00000", 
           "11111", "10010", "11111", "11111", "11111", 
           "11111", "01010", "11111", "11111", "10010", 
           "10010", "11111", "10011", "00001", "00000", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "01010", "10010", "10010", "11111", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "10010", "10010", "10010", "10010", 
           "10010", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "10010", "11111", "11111", "11111", 
           "10010", "01010", "10010", "10010", "10010", 
           "10010", "10010", "11111", "00001", "00000", 
           "11111", "10010", "10010", "10010", "10010", 
           "10010", "01010", "11111", "11111", "11111", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "01010", "10010", "10010", "10010", 
           "10010", "10010", "10011", "00001", "00000", 
           "11111", "10010", "10010", "10010", "10010", 
           "10010", "01010", "11111", "10010", "11111", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "11111", "11111", "11111", "11111", 
           "10010", "01010", "11111", "11111", "10010", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "10010", "10010", "10010", "10010", 
           "10010", "01010", "11111", "11111", "11111", 
           "10010", "11111", "11111", "00001", "00000", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "10010", "10010", "10010", 
           "10010", "10010", "10011", "00001", "00000", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "00001", "00000", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "00001", "00000", 
           "01001", "01001", "01001", "01001", "01001", 
           "01001", "01001", "01001", "01001", "01001", 
           "01001", "01001", "01001", "00001", "00000", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111", 
           "11111", "11111", "11111", "11111", "11111");

	signal query_help : unsigned(4 downto 0);
	signal data_main : std_logic_vector(4 downto 0);
	signal data_win : std_logic_vector(4 downto 0);

begin
    process(clk)
    begin
        if rising_edge(clk) then
            data_main <= pictMem(to_integer(addr));
            data_win <= you_win(to_integer(addr));
            query_help <= unsigned(pictMem(to_integer(query_addr)));
        end if;
    end process;

    query_result <= '0' when query_help > 15 else '1';

	with level_choice select data_out <=
		data_main when '0',
		data_win when others;

end Behavioral;
